module InstructionMemoryCache(
  input         clock,
  input         reset,
  input         io_fetch_0_address_valid,
  input  [63:0] io_fetch_0_address_bits,
  output        io_fetch_0_output_valid,
  output [31:0] io_fetch_0_output_bits,
  input         io_memory_request_ready,
  output        io_memory_request_valid,
  output [63:0] io_memory_request_bits_address,
  input         io_memory_response_valid,
  input  [63:0] io_memory_response_bits_inner
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [63:0] _RAND_42;
  reg [63:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
`endif // RANDOMIZE_REG_INIT
  reg  buf_0_valid; // @[InstructionMemoryCache.scala 41:28]
  reg [59:0] buf_0_upper; // @[InstructionMemoryCache.scala 41:28]
  reg [15:0] buf_0_data_0; // @[InstructionMemoryCache.scala 41:28]
  reg [15:0] buf_0_data_1; // @[InstructionMemoryCache.scala 41:28]
  reg [15:0] buf_0_data_2; // @[InstructionMemoryCache.scala 41:28]
  reg [15:0] buf_0_data_3; // @[InstructionMemoryCache.scala 41:28]
  reg [15:0] buf_0_data_4; // @[InstructionMemoryCache.scala 41:28]
  reg [15:0] buf_0_data_5; // @[InstructionMemoryCache.scala 41:28]
  reg [15:0] buf_0_data_6; // @[InstructionMemoryCache.scala 41:28]
  reg [15:0] buf_0_data_7; // @[InstructionMemoryCache.scala 41:28]
  reg  buf_1_valid; // @[InstructionMemoryCache.scala 41:28]
  reg [59:0] buf_1_upper; // @[InstructionMemoryCache.scala 41:28]
  reg [15:0] buf_1_data_0; // @[InstructionMemoryCache.scala 41:28]
  reg [15:0] buf_1_data_1; // @[InstructionMemoryCache.scala 41:28]
  reg [15:0] buf_1_data_2; // @[InstructionMemoryCache.scala 41:28]
  reg [15:0] buf_1_data_3; // @[InstructionMemoryCache.scala 41:28]
  reg [15:0] buf_1_data_4; // @[InstructionMemoryCache.scala 41:28]
  reg [15:0] buf_1_data_5; // @[InstructionMemoryCache.scala 41:28]
  reg [15:0] buf_1_data_6; // @[InstructionMemoryCache.scala 41:28]
  reg [15:0] buf_1_data_7; // @[InstructionMemoryCache.scala 41:28]
  reg  buf_2_valid; // @[InstructionMemoryCache.scala 41:28]
  reg [59:0] buf_2_upper; // @[InstructionMemoryCache.scala 41:28]
  reg [15:0] buf_2_data_0; // @[InstructionMemoryCache.scala 41:28]
  reg [15:0] buf_2_data_1; // @[InstructionMemoryCache.scala 41:28]
  reg [15:0] buf_2_data_2; // @[InstructionMemoryCache.scala 41:28]
  reg [15:0] buf_2_data_3; // @[InstructionMemoryCache.scala 41:28]
  reg [15:0] buf_2_data_4; // @[InstructionMemoryCache.scala 41:28]
  reg [15:0] buf_2_data_5; // @[InstructionMemoryCache.scala 41:28]
  reg [15:0] buf_2_data_6; // @[InstructionMemoryCache.scala 41:28]
  reg [15:0] buf_2_data_7; // @[InstructionMemoryCache.scala 41:28]
  reg  buf_3_valid; // @[InstructionMemoryCache.scala 41:28]
  reg [59:0] buf_3_upper; // @[InstructionMemoryCache.scala 41:28]
  reg [15:0] buf_3_data_0; // @[InstructionMemoryCache.scala 41:28]
  reg [15:0] buf_3_data_1; // @[InstructionMemoryCache.scala 41:28]
  reg [15:0] buf_3_data_2; // @[InstructionMemoryCache.scala 41:28]
  reg [15:0] buf_3_data_3; // @[InstructionMemoryCache.scala 41:28]
  reg [15:0] buf_3_data_4; // @[InstructionMemoryCache.scala 41:28]
  reg [15:0] buf_3_data_5; // @[InstructionMemoryCache.scala 41:28]
  reg [15:0] buf_3_data_6; // @[InstructionMemoryCache.scala 41:28]
  reg [15:0] buf_3_data_7; // @[InstructionMemoryCache.scala 41:28]
  wire [62:0] lowerAddress = io_fetch_0_address_bits[63:1]; // @[InstructionMemoryCache.scala 46:38]
  wire [62:0] upperAddress = lowerAddress + 63'h1; // @[InstructionMemoryCache.scala 47:37]
  wire  _T_4 = buf_0_valid & lowerAddress[62:3] == buf_0_upper; // @[InstructionMemoryCache.scala 54:34]
  wire [15:0] _GEN_1 = 3'h1 == lowerAddress[2:0] ? buf_0_data_1 : buf_0_data_0; // @[InstructionMemoryCache.scala 55:{19,19}]
  wire [15:0] _GEN_2 = 3'h2 == lowerAddress[2:0] ? buf_0_data_2 : _GEN_1; // @[InstructionMemoryCache.scala 55:{19,19}]
  wire [15:0] _GEN_3 = 3'h3 == lowerAddress[2:0] ? buf_0_data_3 : _GEN_2; // @[InstructionMemoryCache.scala 55:{19,19}]
  wire [15:0] _GEN_4 = 3'h4 == lowerAddress[2:0] ? buf_0_data_4 : _GEN_3; // @[InstructionMemoryCache.scala 55:{19,19}]
  wire [15:0] _GEN_5 = 3'h5 == lowerAddress[2:0] ? buf_0_data_5 : _GEN_4; // @[InstructionMemoryCache.scala 55:{19,19}]
  wire [15:0] _GEN_6 = 3'h6 == lowerAddress[2:0] ? buf_0_data_6 : _GEN_5; // @[InstructionMemoryCache.scala 55:{19,19}]
  wire [15:0] _GEN_7 = 3'h7 == lowerAddress[2:0] ? buf_0_data_7 : _GEN_6; // @[InstructionMemoryCache.scala 55:{19,19}]
  wire [15:0] _GEN_8 = buf_0_valid & lowerAddress[62:3] == buf_0_upper ? _GEN_7 : 16'h0; // @[InstructionMemoryCache.scala 54:70 55:19 48:32]
  wire  _T_12 = lowerAddress[62:3] == buf_1_upper; // @[InstructionMemoryCache.scala 54:57]
  wire [15:0] _GEN_10 = 3'h1 == lowerAddress[2:0] ? buf_1_data_1 : buf_1_data_0; // @[InstructionMemoryCache.scala 55:{19,19}]
  wire [15:0] _GEN_11 = 3'h2 == lowerAddress[2:0] ? buf_1_data_2 : _GEN_10; // @[InstructionMemoryCache.scala 55:{19,19}]
  wire [15:0] _GEN_12 = 3'h3 == lowerAddress[2:0] ? buf_1_data_3 : _GEN_11; // @[InstructionMemoryCache.scala 55:{19,19}]
  wire [15:0] _GEN_13 = 3'h4 == lowerAddress[2:0] ? buf_1_data_4 : _GEN_12; // @[InstructionMemoryCache.scala 55:{19,19}]
  wire [15:0] _GEN_14 = 3'h5 == lowerAddress[2:0] ? buf_1_data_5 : _GEN_13; // @[InstructionMemoryCache.scala 55:{19,19}]
  wire [15:0] _GEN_15 = 3'h6 == lowerAddress[2:0] ? buf_1_data_6 : _GEN_14; // @[InstructionMemoryCache.scala 55:{19,19}]
  wire [15:0] _GEN_16 = 3'h7 == lowerAddress[2:0] ? buf_1_data_7 : _GEN_15; // @[InstructionMemoryCache.scala 55:{19,19}]
  wire [15:0] _GEN_17 = ~(buf_0_valid & lowerAddress[62:3] == buf_0_upper) & buf_1_valid & lowerAddress[62:3] ==
    buf_1_upper ? _GEN_16 : _GEN_8; // @[InstructionMemoryCache.scala 54:70 55:19]
  wire  _T_17 = _T_4 | buf_1_valid & _T_12; // @[InstructionMemoryCache.scala 57:29]
  wire  _T_21 = lowerAddress[62:3] == buf_2_upper; // @[InstructionMemoryCache.scala 54:57]
  wire [15:0] _GEN_19 = 3'h1 == lowerAddress[2:0] ? buf_2_data_1 : buf_2_data_0; // @[InstructionMemoryCache.scala 55:{19,19}]
  wire [15:0] _GEN_20 = 3'h2 == lowerAddress[2:0] ? buf_2_data_2 : _GEN_19; // @[InstructionMemoryCache.scala 55:{19,19}]
  wire [15:0] _GEN_21 = 3'h3 == lowerAddress[2:0] ? buf_2_data_3 : _GEN_20; // @[InstructionMemoryCache.scala 55:{19,19}]
  wire [15:0] _GEN_22 = 3'h4 == lowerAddress[2:0] ? buf_2_data_4 : _GEN_21; // @[InstructionMemoryCache.scala 55:{19,19}]
  wire [15:0] _GEN_23 = 3'h5 == lowerAddress[2:0] ? buf_2_data_5 : _GEN_22; // @[InstructionMemoryCache.scala 55:{19,19}]
  wire [15:0] _GEN_24 = 3'h6 == lowerAddress[2:0] ? buf_2_data_6 : _GEN_23; // @[InstructionMemoryCache.scala 55:{19,19}]
  wire [15:0] _GEN_25 = 3'h7 == lowerAddress[2:0] ? buf_2_data_7 : _GEN_24; // @[InstructionMemoryCache.scala 55:{19,19}]
  wire [15:0] _GEN_26 = ~_T_17 & buf_2_valid & lowerAddress[62:3] == buf_2_upper ? _GEN_25 : _GEN_17; // @[InstructionMemoryCache.scala 54:70 55:19]
  wire  _T_26 = _T_4 | buf_1_valid & _T_12 | buf_2_valid & _T_21; // @[InstructionMemoryCache.scala 57:29]
  wire  _T_30 = lowerAddress[62:3] == buf_3_upper; // @[InstructionMemoryCache.scala 54:57]
  wire [15:0] _GEN_28 = 3'h1 == lowerAddress[2:0] ? buf_3_data_1 : buf_3_data_0; // @[InstructionMemoryCache.scala 55:{19,19}]
  wire [15:0] _GEN_29 = 3'h2 == lowerAddress[2:0] ? buf_3_data_2 : _GEN_28; // @[InstructionMemoryCache.scala 55:{19,19}]
  wire [15:0] _GEN_30 = 3'h3 == lowerAddress[2:0] ? buf_3_data_3 : _GEN_29; // @[InstructionMemoryCache.scala 55:{19,19}]
  wire [15:0] _GEN_31 = 3'h4 == lowerAddress[2:0] ? buf_3_data_4 : _GEN_30; // @[InstructionMemoryCache.scala 55:{19,19}]
  wire [15:0] _GEN_32 = 3'h5 == lowerAddress[2:0] ? buf_3_data_5 : _GEN_31; // @[InstructionMemoryCache.scala 55:{19,19}]
  wire [15:0] _GEN_33 = 3'h6 == lowerAddress[2:0] ? buf_3_data_6 : _GEN_32; // @[InstructionMemoryCache.scala 55:{19,19}]
  wire [15:0] _GEN_34 = 3'h7 == lowerAddress[2:0] ? buf_3_data_7 : _GEN_33; // @[InstructionMemoryCache.scala 55:{19,19}]
  wire [15:0] lowerData = ~_T_26 & buf_3_valid & lowerAddress[62:3] == buf_3_upper ? _GEN_34 : _GEN_26; // @[InstructionMemoryCache.scala 54:70 55:19]
  wire  _T_35 = _T_4 | buf_1_valid & _T_12 | buf_2_valid & _T_21 | buf_3_valid & _T_30; // @[InstructionMemoryCache.scala 57:29]
  wire  _T_40 = buf_0_valid & upperAddress[62:3] == buf_0_upper; // @[InstructionMemoryCache.scala 62:35]
  wire [15:0] _GEN_37 = 3'h1 == upperAddress[2:0] ? buf_0_data_1 : buf_0_data_0; // @[InstructionMemoryCache.scala 63:{19,19}]
  wire [15:0] _GEN_38 = 3'h2 == upperAddress[2:0] ? buf_0_data_2 : _GEN_37; // @[InstructionMemoryCache.scala 63:{19,19}]
  wire [15:0] _GEN_39 = 3'h3 == upperAddress[2:0] ? buf_0_data_3 : _GEN_38; // @[InstructionMemoryCache.scala 63:{19,19}]
  wire [15:0] _GEN_40 = 3'h4 == upperAddress[2:0] ? buf_0_data_4 : _GEN_39; // @[InstructionMemoryCache.scala 63:{19,19}]
  wire [15:0] _GEN_41 = 3'h5 == upperAddress[2:0] ? buf_0_data_5 : _GEN_40; // @[InstructionMemoryCache.scala 63:{19,19}]
  wire [15:0] _GEN_42 = 3'h6 == upperAddress[2:0] ? buf_0_data_6 : _GEN_41; // @[InstructionMemoryCache.scala 63:{19,19}]
  wire [15:0] _GEN_43 = 3'h7 == upperAddress[2:0] ? buf_0_data_7 : _GEN_42; // @[InstructionMemoryCache.scala 63:{19,19}]
  wire [15:0] _GEN_44 = buf_0_valid & upperAddress[62:3] == buf_0_upper ? _GEN_43 : 16'h0; // @[InstructionMemoryCache.scala 62:71 63:19 49:32]
  wire  _T_48 = upperAddress[62:3] == buf_1_upper; // @[InstructionMemoryCache.scala 62:58]
  wire [15:0] _GEN_46 = 3'h1 == upperAddress[2:0] ? buf_1_data_1 : buf_1_data_0; // @[InstructionMemoryCache.scala 63:{19,19}]
  wire [15:0] _GEN_47 = 3'h2 == upperAddress[2:0] ? buf_1_data_2 : _GEN_46; // @[InstructionMemoryCache.scala 63:{19,19}]
  wire [15:0] _GEN_48 = 3'h3 == upperAddress[2:0] ? buf_1_data_3 : _GEN_47; // @[InstructionMemoryCache.scala 63:{19,19}]
  wire [15:0] _GEN_49 = 3'h4 == upperAddress[2:0] ? buf_1_data_4 : _GEN_48; // @[InstructionMemoryCache.scala 63:{19,19}]
  wire [15:0] _GEN_50 = 3'h5 == upperAddress[2:0] ? buf_1_data_5 : _GEN_49; // @[InstructionMemoryCache.scala 63:{19,19}]
  wire [15:0] _GEN_51 = 3'h6 == upperAddress[2:0] ? buf_1_data_6 : _GEN_50; // @[InstructionMemoryCache.scala 63:{19,19}]
  wire [15:0] _GEN_52 = 3'h7 == upperAddress[2:0] ? buf_1_data_7 : _GEN_51; // @[InstructionMemoryCache.scala 63:{19,19}]
  wire [15:0] _GEN_53 = ~(buf_0_valid & upperAddress[62:3] == buf_0_upper) & buf_1_valid & upperAddress[62:3] ==
    buf_1_upper ? _GEN_52 : _GEN_44; // @[InstructionMemoryCache.scala 62:71 63:19]
  wire  _T_53 = _T_40 | buf_1_valid & _T_48; // @[InstructionMemoryCache.scala 65:31]
  wire  _T_57 = upperAddress[62:3] == buf_2_upper; // @[InstructionMemoryCache.scala 62:58]
  wire [15:0] _GEN_55 = 3'h1 == upperAddress[2:0] ? buf_2_data_1 : buf_2_data_0; // @[InstructionMemoryCache.scala 63:{19,19}]
  wire [15:0] _GEN_56 = 3'h2 == upperAddress[2:0] ? buf_2_data_2 : _GEN_55; // @[InstructionMemoryCache.scala 63:{19,19}]
  wire [15:0] _GEN_57 = 3'h3 == upperAddress[2:0] ? buf_2_data_3 : _GEN_56; // @[InstructionMemoryCache.scala 63:{19,19}]
  wire [15:0] _GEN_58 = 3'h4 == upperAddress[2:0] ? buf_2_data_4 : _GEN_57; // @[InstructionMemoryCache.scala 63:{19,19}]
  wire [15:0] _GEN_59 = 3'h5 == upperAddress[2:0] ? buf_2_data_5 : _GEN_58; // @[InstructionMemoryCache.scala 63:{19,19}]
  wire [15:0] _GEN_60 = 3'h6 == upperAddress[2:0] ? buf_2_data_6 : _GEN_59; // @[InstructionMemoryCache.scala 63:{19,19}]
  wire [15:0] _GEN_61 = 3'h7 == upperAddress[2:0] ? buf_2_data_7 : _GEN_60; // @[InstructionMemoryCache.scala 63:{19,19}]
  wire [15:0] _GEN_62 = ~_T_53 & buf_2_valid & upperAddress[62:3] == buf_2_upper ? _GEN_61 : _GEN_53; // @[InstructionMemoryCache.scala 62:71 63:19]
  wire  _T_62 = _T_40 | buf_1_valid & _T_48 | buf_2_valid & _T_57; // @[InstructionMemoryCache.scala 65:31]
  wire  _T_66 = upperAddress[62:3] == buf_3_upper; // @[InstructionMemoryCache.scala 62:58]
  wire [15:0] _GEN_64 = 3'h1 == upperAddress[2:0] ? buf_3_data_1 : buf_3_data_0; // @[InstructionMemoryCache.scala 63:{19,19}]
  wire [15:0] _GEN_65 = 3'h2 == upperAddress[2:0] ? buf_3_data_2 : _GEN_64; // @[InstructionMemoryCache.scala 63:{19,19}]
  wire [15:0] _GEN_66 = 3'h3 == upperAddress[2:0] ? buf_3_data_3 : _GEN_65; // @[InstructionMemoryCache.scala 63:{19,19}]
  wire [15:0] _GEN_67 = 3'h4 == upperAddress[2:0] ? buf_3_data_4 : _GEN_66; // @[InstructionMemoryCache.scala 63:{19,19}]
  wire [15:0] _GEN_68 = 3'h5 == upperAddress[2:0] ? buf_3_data_5 : _GEN_67; // @[InstructionMemoryCache.scala 63:{19,19}]
  wire [15:0] _GEN_69 = 3'h6 == upperAddress[2:0] ? buf_3_data_6 : _GEN_68; // @[InstructionMemoryCache.scala 63:{19,19}]
  wire [15:0] _GEN_70 = 3'h7 == upperAddress[2:0] ? buf_3_data_7 : _GEN_69; // @[InstructionMemoryCache.scala 63:{19,19}]
  wire [15:0] upperData = ~_T_62 & buf_3_valid & upperAddress[62:3] == buf_3_upper ? _GEN_70 : _GEN_62; // @[InstructionMemoryCache.scala 62:71 63:19]
  wire  _T_71 = _T_40 | buf_1_valid & _T_48 | buf_2_valid & _T_57 | buf_3_valid & _T_66; // @[InstructionMemoryCache.scala 65:31]
  wire  _T_72 = ~_T_35; // @[InstructionMemoryCache.scala 72:12]
  wire  _T_75 = ~_T_71; // @[InstructionMemoryCache.scala 74:18]
  wire [59:0] _GEN_72 = ~_T_71 ? upperAddress[62:3] : 60'h0; // @[InstructionMemoryCache.scala 74:46 75:17 43:36]
  wire [59:0] _GEN_73 = ~_T_35 ? lowerAddress[62:3] : _GEN_72; // @[InstructionMemoryCache.scala 72:39 73:17]
  wire [59:0] request = io_fetch_0_address_valid ? _GEN_73 : 60'h0; // @[InstructionMemoryCache.scala 71:27 43:36]
  wire  _T_81 = (_T_72 | _T_75) & io_fetch_0_address_valid; // @[InstructionMemoryCache.scala 78:60]
  reg  state; // @[InstructionMemoryCache.scala 82:30]
  reg  readIndex; // @[InstructionMemoryCache.scala 83:30]
  reg [59:0] requested; // @[InstructionMemoryCache.scala 84:34]
  reg [63:0] transaction_address; // @[InstructionMemoryCache.scala 85:32]
  reg  requestDone; // @[InstructionMemoryCache.scala 86:32]
  wire [63:0] tmp_transaction_address = {request,4'h0}; // @[Cat.scala 33:92]
  wire  _GEN_75 = _T_81 & ~state | state; // @[InstructionMemoryCache.scala 88:41 89:11 82:30]
  wire  _GEN_77 = _T_81 & ~state ? 1'h0 : readIndex; // @[InstructionMemoryCache.scala 88:41 91:15 83:30]
  wire  _GEN_85 = _T_81 & ~state ? 1'h0 : requestDone; // @[InstructionMemoryCache.scala 88:41 99:17 86:32]
  reg [1:0] head; // @[InstructionMemoryCache.scala 104:29]
  wire  _T_86 = ~requestDone; // @[InstructionMemoryCache.scala 106:10]
  wire  _GEN_86 = io_memory_request_ready | _GEN_85; // @[InstructionMemoryCache.scala 109:37 110:21]
  wire  _GEN_96 = 2'h0 == head ? 1'h0 : buf_0_valid; // @[InstructionMemoryCache.scala 115:{23,23} 41:28]
  wire  _GEN_97 = 2'h1 == head ? 1'h0 : buf_1_valid; // @[InstructionMemoryCache.scala 115:{23,23} 41:28]
  wire  _GEN_98 = 2'h2 == head ? 1'h0 : buf_2_valid; // @[InstructionMemoryCache.scala 115:{23,23} 41:28]
  wire  _GEN_99 = 2'h3 == head ? 1'h0 : buf_3_valid; // @[InstructionMemoryCache.scala 115:{23,23} 41:28]
  wire [2:0] _T_87 = {readIndex,2'h0}; // @[InstructionMemoryCache.scala 117:34]
  wire  _GEN_341 = 2'h0 == head; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [15:0] _GEN_100 = 2'h0 == head & 3'h0 == _T_87 ? io_memory_response_bits_inner[15:0] : buf_0_data_0; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [15:0] _GEN_101 = 2'h0 == head & 3'h1 == _T_87 ? io_memory_response_bits_inner[15:0] : buf_0_data_1; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [15:0] _GEN_102 = 2'h0 == head & 3'h2 == _T_87 ? io_memory_response_bits_inner[15:0] : buf_0_data_2; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [15:0] _GEN_103 = 2'h0 == head & 3'h3 == _T_87 ? io_memory_response_bits_inner[15:0] : buf_0_data_3; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [15:0] _GEN_104 = 2'h0 == head & 3'h4 == _T_87 ? io_memory_response_bits_inner[15:0] : buf_0_data_4; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [15:0] _GEN_105 = 2'h0 == head & 3'h5 == _T_87 ? io_memory_response_bits_inner[15:0] : buf_0_data_5; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [15:0] _GEN_106 = 2'h0 == head & 3'h6 == _T_87 ? io_memory_response_bits_inner[15:0] : buf_0_data_6; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [15:0] _GEN_107 = 2'h0 == head & 3'h7 == _T_87 ? io_memory_response_bits_inner[15:0] : buf_0_data_7; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire  _GEN_357 = 2'h1 == head; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [15:0] _GEN_108 = 2'h1 == head & 3'h0 == _T_87 ? io_memory_response_bits_inner[15:0] : buf_1_data_0; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [15:0] _GEN_109 = 2'h1 == head & 3'h1 == _T_87 ? io_memory_response_bits_inner[15:0] : buf_1_data_1; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [15:0] _GEN_110 = 2'h1 == head & 3'h2 == _T_87 ? io_memory_response_bits_inner[15:0] : buf_1_data_2; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [15:0] _GEN_111 = 2'h1 == head & 3'h3 == _T_87 ? io_memory_response_bits_inner[15:0] : buf_1_data_3; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [15:0] _GEN_112 = 2'h1 == head & 3'h4 == _T_87 ? io_memory_response_bits_inner[15:0] : buf_1_data_4; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [15:0] _GEN_113 = 2'h1 == head & 3'h5 == _T_87 ? io_memory_response_bits_inner[15:0] : buf_1_data_5; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [15:0] _GEN_114 = 2'h1 == head & 3'h6 == _T_87 ? io_memory_response_bits_inner[15:0] : buf_1_data_6; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [15:0] _GEN_115 = 2'h1 == head & 3'h7 == _T_87 ? io_memory_response_bits_inner[15:0] : buf_1_data_7; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire  _GEN_373 = 2'h2 == head; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [15:0] _GEN_116 = 2'h2 == head & 3'h0 == _T_87 ? io_memory_response_bits_inner[15:0] : buf_2_data_0; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [15:0] _GEN_117 = 2'h2 == head & 3'h1 == _T_87 ? io_memory_response_bits_inner[15:0] : buf_2_data_1; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [15:0] _GEN_118 = 2'h2 == head & 3'h2 == _T_87 ? io_memory_response_bits_inner[15:0] : buf_2_data_2; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [15:0] _GEN_119 = 2'h2 == head & 3'h3 == _T_87 ? io_memory_response_bits_inner[15:0] : buf_2_data_3; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [15:0] _GEN_120 = 2'h2 == head & 3'h4 == _T_87 ? io_memory_response_bits_inner[15:0] : buf_2_data_4; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [15:0] _GEN_121 = 2'h2 == head & 3'h5 == _T_87 ? io_memory_response_bits_inner[15:0] : buf_2_data_5; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [15:0] _GEN_122 = 2'h2 == head & 3'h6 == _T_87 ? io_memory_response_bits_inner[15:0] : buf_2_data_6; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [15:0] _GEN_123 = 2'h2 == head & 3'h7 == _T_87 ? io_memory_response_bits_inner[15:0] : buf_2_data_7; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire  _GEN_389 = 2'h3 == head; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [15:0] _GEN_124 = 2'h3 == head & 3'h0 == _T_87 ? io_memory_response_bits_inner[15:0] : buf_3_data_0; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [15:0] _GEN_125 = 2'h3 == head & 3'h1 == _T_87 ? io_memory_response_bits_inner[15:0] : buf_3_data_1; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [15:0] _GEN_126 = 2'h3 == head & 3'h2 == _T_87 ? io_memory_response_bits_inner[15:0] : buf_3_data_2; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [15:0] _GEN_127 = 2'h3 == head & 3'h3 == _T_87 ? io_memory_response_bits_inner[15:0] : buf_3_data_3; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [15:0] _GEN_128 = 2'h3 == head & 3'h4 == _T_87 ? io_memory_response_bits_inner[15:0] : buf_3_data_4; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [15:0] _GEN_129 = 2'h3 == head & 3'h5 == _T_87 ? io_memory_response_bits_inner[15:0] : buf_3_data_5; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [15:0] _GEN_130 = 2'h3 == head & 3'h6 == _T_87 ? io_memory_response_bits_inner[15:0] : buf_3_data_6; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [15:0] _GEN_131 = 2'h3 == head & 3'h7 == _T_87 ? io_memory_response_bits_inner[15:0] : buf_3_data_7; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [2:0] _T_88 = {readIndex,2'h1}; // @[InstructionMemoryCache.scala 117:34]
  wire [15:0] _GEN_132 = _GEN_341 & 3'h0 == _T_88 ? io_memory_response_bits_inner[31:16] : _GEN_100; // @[InstructionMemoryCache.scala 117:{47,47}]
  wire [15:0] _GEN_133 = _GEN_341 & 3'h1 == _T_88 ? io_memory_response_bits_inner[31:16] : _GEN_101; // @[InstructionMemoryCache.scala 117:{47,47}]
  wire [15:0] _GEN_134 = _GEN_341 & 3'h2 == _T_88 ? io_memory_response_bits_inner[31:16] : _GEN_102; // @[InstructionMemoryCache.scala 117:{47,47}]
  wire [15:0] _GEN_135 = _GEN_341 & 3'h3 == _T_88 ? io_memory_response_bits_inner[31:16] : _GEN_103; // @[InstructionMemoryCache.scala 117:{47,47}]
  wire [15:0] _GEN_136 = _GEN_341 & 3'h4 == _T_88 ? io_memory_response_bits_inner[31:16] : _GEN_104; // @[InstructionMemoryCache.scala 117:{47,47}]
  wire [15:0] _GEN_137 = _GEN_341 & 3'h5 == _T_88 ? io_memory_response_bits_inner[31:16] : _GEN_105; // @[InstructionMemoryCache.scala 117:{47,47}]
  wire [15:0] _GEN_138 = _GEN_341 & 3'h6 == _T_88 ? io_memory_response_bits_inner[31:16] : _GEN_106; // @[InstructionMemoryCache.scala 117:{47,47}]
  wire [15:0] _GEN_139 = _GEN_341 & 3'h7 == _T_88 ? io_memory_response_bits_inner[31:16] : _GEN_107; // @[InstructionMemoryCache.scala 117:{47,47}]
  wire [15:0] _GEN_140 = _GEN_357 & 3'h0 == _T_88 ? io_memory_response_bits_inner[31:16] : _GEN_108; // @[InstructionMemoryCache.scala 117:{47,47}]
  wire [15:0] _GEN_141 = _GEN_357 & 3'h1 == _T_88 ? io_memory_response_bits_inner[31:16] : _GEN_109; // @[InstructionMemoryCache.scala 117:{47,47}]
  wire [15:0] _GEN_142 = _GEN_357 & 3'h2 == _T_88 ? io_memory_response_bits_inner[31:16] : _GEN_110; // @[InstructionMemoryCache.scala 117:{47,47}]
  wire [15:0] _GEN_143 = _GEN_357 & 3'h3 == _T_88 ? io_memory_response_bits_inner[31:16] : _GEN_111; // @[InstructionMemoryCache.scala 117:{47,47}]
  wire [15:0] _GEN_144 = _GEN_357 & 3'h4 == _T_88 ? io_memory_response_bits_inner[31:16] : _GEN_112; // @[InstructionMemoryCache.scala 117:{47,47}]
  wire [15:0] _GEN_145 = _GEN_357 & 3'h5 == _T_88 ? io_memory_response_bits_inner[31:16] : _GEN_113; // @[InstructionMemoryCache.scala 117:{47,47}]
  wire [15:0] _GEN_146 = _GEN_357 & 3'h6 == _T_88 ? io_memory_response_bits_inner[31:16] : _GEN_114; // @[InstructionMemoryCache.scala 117:{47,47}]
  wire [15:0] _GEN_147 = _GEN_357 & 3'h7 == _T_88 ? io_memory_response_bits_inner[31:16] : _GEN_115; // @[InstructionMemoryCache.scala 117:{47,47}]
  wire [15:0] _GEN_148 = _GEN_373 & 3'h0 == _T_88 ? io_memory_response_bits_inner[31:16] : _GEN_116; // @[InstructionMemoryCache.scala 117:{47,47}]
  wire [15:0] _GEN_149 = _GEN_373 & 3'h1 == _T_88 ? io_memory_response_bits_inner[31:16] : _GEN_117; // @[InstructionMemoryCache.scala 117:{47,47}]
  wire [15:0] _GEN_150 = _GEN_373 & 3'h2 == _T_88 ? io_memory_response_bits_inner[31:16] : _GEN_118; // @[InstructionMemoryCache.scala 117:{47,47}]
  wire [15:0] _GEN_151 = _GEN_373 & 3'h3 == _T_88 ? io_memory_response_bits_inner[31:16] : _GEN_119; // @[InstructionMemoryCache.scala 117:{47,47}]
  wire [15:0] _GEN_152 = _GEN_373 & 3'h4 == _T_88 ? io_memory_response_bits_inner[31:16] : _GEN_120; // @[InstructionMemoryCache.scala 117:{47,47}]
  wire [15:0] _GEN_153 = _GEN_373 & 3'h5 == _T_88 ? io_memory_response_bits_inner[31:16] : _GEN_121; // @[InstructionMemoryCache.scala 117:{47,47}]
  wire [15:0] _GEN_154 = _GEN_373 & 3'h6 == _T_88 ? io_memory_response_bits_inner[31:16] : _GEN_122; // @[InstructionMemoryCache.scala 117:{47,47}]
  wire [15:0] _GEN_155 = _GEN_373 & 3'h7 == _T_88 ? io_memory_response_bits_inner[31:16] : _GEN_123; // @[InstructionMemoryCache.scala 117:{47,47}]
  wire [15:0] _GEN_156 = _GEN_389 & 3'h0 == _T_88 ? io_memory_response_bits_inner[31:16] : _GEN_124; // @[InstructionMemoryCache.scala 117:{47,47}]
  wire [15:0] _GEN_157 = _GEN_389 & 3'h1 == _T_88 ? io_memory_response_bits_inner[31:16] : _GEN_125; // @[InstructionMemoryCache.scala 117:{47,47}]
  wire [15:0] _GEN_158 = _GEN_389 & 3'h2 == _T_88 ? io_memory_response_bits_inner[31:16] : _GEN_126; // @[InstructionMemoryCache.scala 117:{47,47}]
  wire [15:0] _GEN_159 = _GEN_389 & 3'h3 == _T_88 ? io_memory_response_bits_inner[31:16] : _GEN_127; // @[InstructionMemoryCache.scala 117:{47,47}]
  wire [15:0] _GEN_160 = _GEN_389 & 3'h4 == _T_88 ? io_memory_response_bits_inner[31:16] : _GEN_128; // @[InstructionMemoryCache.scala 117:{47,47}]
  wire [15:0] _GEN_161 = _GEN_389 & 3'h5 == _T_88 ? io_memory_response_bits_inner[31:16] : _GEN_129; // @[InstructionMemoryCache.scala 117:{47,47}]
  wire [15:0] _GEN_162 = _GEN_389 & 3'h6 == _T_88 ? io_memory_response_bits_inner[31:16] : _GEN_130; // @[InstructionMemoryCache.scala 117:{47,47}]
  wire [15:0] _GEN_163 = _GEN_389 & 3'h7 == _T_88 ? io_memory_response_bits_inner[31:16] : _GEN_131; // @[InstructionMemoryCache.scala 117:{47,47}]
  wire [2:0] _T_89 = {readIndex,2'h2}; // @[InstructionMemoryCache.scala 117:34]
  wire [2:0] _T_90 = {readIndex,2'h3}; // @[InstructionMemoryCache.scala 117:34]
  wire  _GEN_228 = _GEN_341 | _GEN_96; // @[InstructionMemoryCache.scala 123:{25,25}]
  wire  _GEN_229 = _GEN_357 | _GEN_97; // @[InstructionMemoryCache.scala 123:{25,25}]
  wire  _GEN_230 = _GEN_373 | _GEN_98; // @[InstructionMemoryCache.scala 123:{25,25}]
  wire  _GEN_231 = _GEN_389 | _GEN_99; // @[InstructionMemoryCache.scala 123:{25,25}]
  wire [1:0] _head_T_1 = head + 2'h1; // @[InstructionMemoryCache.scala 125:22]
  assign io_fetch_0_output_valid = _T_35 & _T_71; // @[InstructionMemoryCache.scala 68:33]
  assign io_fetch_0_output_bits = {upperData,lowerData}; // @[InstructionMemoryCache.scala 69:32]
  assign io_memory_request_valid = state & _T_86; // @[InstructionMemoryCache.scala 102:27 105:30]
  assign io_memory_request_bits_address = transaction_address; // @[InstructionMemoryCache.scala 106:24 108:30]
  always @(posedge clock) begin
    if (reset) begin // @[InstructionMemoryCache.scala 41:28]
      buf_0_valid <= 1'h0; // @[InstructionMemoryCache.scala 41:28]
    end else if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (readIndex) begin // @[InstructionMemoryCache.scala 121:31]
          buf_0_valid <= _GEN_228;
        end else begin
          buf_0_valid <= _GEN_96;
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (readIndex) begin // @[InstructionMemoryCache.scala 121:31]
          if (2'h0 == head) begin // @[InstructionMemoryCache.scala 124:25]
            buf_0_upper <= requested; // @[InstructionMemoryCache.scala 124:25]
          end
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (_GEN_341 & 3'h0 == _T_90) begin // @[InstructionMemoryCache.scala 117:47]
          buf_0_data_0 <= io_memory_response_bits_inner[63:48]; // @[InstructionMemoryCache.scala 117:47]
        end else if (_GEN_341 & 3'h0 == _T_89) begin // @[InstructionMemoryCache.scala 117:47]
          buf_0_data_0 <= io_memory_response_bits_inner[47:32]; // @[InstructionMemoryCache.scala 117:47]
        end else begin
          buf_0_data_0 <= _GEN_132;
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (_GEN_341 & 3'h1 == _T_90) begin // @[InstructionMemoryCache.scala 117:47]
          buf_0_data_1 <= io_memory_response_bits_inner[63:48]; // @[InstructionMemoryCache.scala 117:47]
        end else if (_GEN_341 & 3'h1 == _T_89) begin // @[InstructionMemoryCache.scala 117:47]
          buf_0_data_1 <= io_memory_response_bits_inner[47:32]; // @[InstructionMemoryCache.scala 117:47]
        end else begin
          buf_0_data_1 <= _GEN_133;
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (_GEN_341 & 3'h2 == _T_90) begin // @[InstructionMemoryCache.scala 117:47]
          buf_0_data_2 <= io_memory_response_bits_inner[63:48]; // @[InstructionMemoryCache.scala 117:47]
        end else if (_GEN_341 & 3'h2 == _T_89) begin // @[InstructionMemoryCache.scala 117:47]
          buf_0_data_2 <= io_memory_response_bits_inner[47:32]; // @[InstructionMemoryCache.scala 117:47]
        end else begin
          buf_0_data_2 <= _GEN_134;
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (_GEN_341 & 3'h3 == _T_90) begin // @[InstructionMemoryCache.scala 117:47]
          buf_0_data_3 <= io_memory_response_bits_inner[63:48]; // @[InstructionMemoryCache.scala 117:47]
        end else if (_GEN_341 & 3'h3 == _T_89) begin // @[InstructionMemoryCache.scala 117:47]
          buf_0_data_3 <= io_memory_response_bits_inner[47:32]; // @[InstructionMemoryCache.scala 117:47]
        end else begin
          buf_0_data_3 <= _GEN_135;
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (_GEN_341 & 3'h4 == _T_90) begin // @[InstructionMemoryCache.scala 117:47]
          buf_0_data_4 <= io_memory_response_bits_inner[63:48]; // @[InstructionMemoryCache.scala 117:47]
        end else if (_GEN_341 & 3'h4 == _T_89) begin // @[InstructionMemoryCache.scala 117:47]
          buf_0_data_4 <= io_memory_response_bits_inner[47:32]; // @[InstructionMemoryCache.scala 117:47]
        end else begin
          buf_0_data_4 <= _GEN_136;
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (_GEN_341 & 3'h5 == _T_90) begin // @[InstructionMemoryCache.scala 117:47]
          buf_0_data_5 <= io_memory_response_bits_inner[63:48]; // @[InstructionMemoryCache.scala 117:47]
        end else if (_GEN_341 & 3'h5 == _T_89) begin // @[InstructionMemoryCache.scala 117:47]
          buf_0_data_5 <= io_memory_response_bits_inner[47:32]; // @[InstructionMemoryCache.scala 117:47]
        end else begin
          buf_0_data_5 <= _GEN_137;
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (_GEN_341 & 3'h6 == _T_90) begin // @[InstructionMemoryCache.scala 117:47]
          buf_0_data_6 <= io_memory_response_bits_inner[63:48]; // @[InstructionMemoryCache.scala 117:47]
        end else if (_GEN_341 & 3'h6 == _T_89) begin // @[InstructionMemoryCache.scala 117:47]
          buf_0_data_6 <= io_memory_response_bits_inner[47:32]; // @[InstructionMemoryCache.scala 117:47]
        end else begin
          buf_0_data_6 <= _GEN_138;
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (_GEN_341 & 3'h7 == _T_90) begin // @[InstructionMemoryCache.scala 117:47]
          buf_0_data_7 <= io_memory_response_bits_inner[63:48]; // @[InstructionMemoryCache.scala 117:47]
        end else if (_GEN_341 & 3'h7 == _T_89) begin // @[InstructionMemoryCache.scala 117:47]
          buf_0_data_7 <= io_memory_response_bits_inner[47:32]; // @[InstructionMemoryCache.scala 117:47]
        end else begin
          buf_0_data_7 <= _GEN_139;
        end
      end
    end
    if (reset) begin // @[InstructionMemoryCache.scala 41:28]
      buf_1_valid <= 1'h0; // @[InstructionMemoryCache.scala 41:28]
    end else if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (readIndex) begin // @[InstructionMemoryCache.scala 121:31]
          buf_1_valid <= _GEN_229;
        end else begin
          buf_1_valid <= _GEN_97;
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (readIndex) begin // @[InstructionMemoryCache.scala 121:31]
          if (2'h1 == head) begin // @[InstructionMemoryCache.scala 124:25]
            buf_1_upper <= requested; // @[InstructionMemoryCache.scala 124:25]
          end
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (_GEN_357 & 3'h0 == _T_90) begin // @[InstructionMemoryCache.scala 117:47]
          buf_1_data_0 <= io_memory_response_bits_inner[63:48]; // @[InstructionMemoryCache.scala 117:47]
        end else if (_GEN_357 & 3'h0 == _T_89) begin // @[InstructionMemoryCache.scala 117:47]
          buf_1_data_0 <= io_memory_response_bits_inner[47:32]; // @[InstructionMemoryCache.scala 117:47]
        end else begin
          buf_1_data_0 <= _GEN_140;
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (_GEN_357 & 3'h1 == _T_90) begin // @[InstructionMemoryCache.scala 117:47]
          buf_1_data_1 <= io_memory_response_bits_inner[63:48]; // @[InstructionMemoryCache.scala 117:47]
        end else if (_GEN_357 & 3'h1 == _T_89) begin // @[InstructionMemoryCache.scala 117:47]
          buf_1_data_1 <= io_memory_response_bits_inner[47:32]; // @[InstructionMemoryCache.scala 117:47]
        end else begin
          buf_1_data_1 <= _GEN_141;
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (_GEN_357 & 3'h2 == _T_90) begin // @[InstructionMemoryCache.scala 117:47]
          buf_1_data_2 <= io_memory_response_bits_inner[63:48]; // @[InstructionMemoryCache.scala 117:47]
        end else if (_GEN_357 & 3'h2 == _T_89) begin // @[InstructionMemoryCache.scala 117:47]
          buf_1_data_2 <= io_memory_response_bits_inner[47:32]; // @[InstructionMemoryCache.scala 117:47]
        end else begin
          buf_1_data_2 <= _GEN_142;
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (_GEN_357 & 3'h3 == _T_90) begin // @[InstructionMemoryCache.scala 117:47]
          buf_1_data_3 <= io_memory_response_bits_inner[63:48]; // @[InstructionMemoryCache.scala 117:47]
        end else if (_GEN_357 & 3'h3 == _T_89) begin // @[InstructionMemoryCache.scala 117:47]
          buf_1_data_3 <= io_memory_response_bits_inner[47:32]; // @[InstructionMemoryCache.scala 117:47]
        end else begin
          buf_1_data_3 <= _GEN_143;
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (_GEN_357 & 3'h4 == _T_90) begin // @[InstructionMemoryCache.scala 117:47]
          buf_1_data_4 <= io_memory_response_bits_inner[63:48]; // @[InstructionMemoryCache.scala 117:47]
        end else if (_GEN_357 & 3'h4 == _T_89) begin // @[InstructionMemoryCache.scala 117:47]
          buf_1_data_4 <= io_memory_response_bits_inner[47:32]; // @[InstructionMemoryCache.scala 117:47]
        end else begin
          buf_1_data_4 <= _GEN_144;
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (_GEN_357 & 3'h5 == _T_90) begin // @[InstructionMemoryCache.scala 117:47]
          buf_1_data_5 <= io_memory_response_bits_inner[63:48]; // @[InstructionMemoryCache.scala 117:47]
        end else if (_GEN_357 & 3'h5 == _T_89) begin // @[InstructionMemoryCache.scala 117:47]
          buf_1_data_5 <= io_memory_response_bits_inner[47:32]; // @[InstructionMemoryCache.scala 117:47]
        end else begin
          buf_1_data_5 <= _GEN_145;
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (_GEN_357 & 3'h6 == _T_90) begin // @[InstructionMemoryCache.scala 117:47]
          buf_1_data_6 <= io_memory_response_bits_inner[63:48]; // @[InstructionMemoryCache.scala 117:47]
        end else if (_GEN_357 & 3'h6 == _T_89) begin // @[InstructionMemoryCache.scala 117:47]
          buf_1_data_6 <= io_memory_response_bits_inner[47:32]; // @[InstructionMemoryCache.scala 117:47]
        end else begin
          buf_1_data_6 <= _GEN_146;
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (_GEN_357 & 3'h7 == _T_90) begin // @[InstructionMemoryCache.scala 117:47]
          buf_1_data_7 <= io_memory_response_bits_inner[63:48]; // @[InstructionMemoryCache.scala 117:47]
        end else if (_GEN_357 & 3'h7 == _T_89) begin // @[InstructionMemoryCache.scala 117:47]
          buf_1_data_7 <= io_memory_response_bits_inner[47:32]; // @[InstructionMemoryCache.scala 117:47]
        end else begin
          buf_1_data_7 <= _GEN_147;
        end
      end
    end
    if (reset) begin // @[InstructionMemoryCache.scala 41:28]
      buf_2_valid <= 1'h0; // @[InstructionMemoryCache.scala 41:28]
    end else if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (readIndex) begin // @[InstructionMemoryCache.scala 121:31]
          buf_2_valid <= _GEN_230;
        end else begin
          buf_2_valid <= _GEN_98;
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (readIndex) begin // @[InstructionMemoryCache.scala 121:31]
          if (2'h2 == head) begin // @[InstructionMemoryCache.scala 124:25]
            buf_2_upper <= requested; // @[InstructionMemoryCache.scala 124:25]
          end
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (_GEN_373 & 3'h0 == _T_90) begin // @[InstructionMemoryCache.scala 117:47]
          buf_2_data_0 <= io_memory_response_bits_inner[63:48]; // @[InstructionMemoryCache.scala 117:47]
        end else if (_GEN_373 & 3'h0 == _T_89) begin // @[InstructionMemoryCache.scala 117:47]
          buf_2_data_0 <= io_memory_response_bits_inner[47:32]; // @[InstructionMemoryCache.scala 117:47]
        end else begin
          buf_2_data_0 <= _GEN_148;
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (_GEN_373 & 3'h1 == _T_90) begin // @[InstructionMemoryCache.scala 117:47]
          buf_2_data_1 <= io_memory_response_bits_inner[63:48]; // @[InstructionMemoryCache.scala 117:47]
        end else if (_GEN_373 & 3'h1 == _T_89) begin // @[InstructionMemoryCache.scala 117:47]
          buf_2_data_1 <= io_memory_response_bits_inner[47:32]; // @[InstructionMemoryCache.scala 117:47]
        end else begin
          buf_2_data_1 <= _GEN_149;
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (_GEN_373 & 3'h2 == _T_90) begin // @[InstructionMemoryCache.scala 117:47]
          buf_2_data_2 <= io_memory_response_bits_inner[63:48]; // @[InstructionMemoryCache.scala 117:47]
        end else if (_GEN_373 & 3'h2 == _T_89) begin // @[InstructionMemoryCache.scala 117:47]
          buf_2_data_2 <= io_memory_response_bits_inner[47:32]; // @[InstructionMemoryCache.scala 117:47]
        end else begin
          buf_2_data_2 <= _GEN_150;
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (_GEN_373 & 3'h3 == _T_90) begin // @[InstructionMemoryCache.scala 117:47]
          buf_2_data_3 <= io_memory_response_bits_inner[63:48]; // @[InstructionMemoryCache.scala 117:47]
        end else if (_GEN_373 & 3'h3 == _T_89) begin // @[InstructionMemoryCache.scala 117:47]
          buf_2_data_3 <= io_memory_response_bits_inner[47:32]; // @[InstructionMemoryCache.scala 117:47]
        end else begin
          buf_2_data_3 <= _GEN_151;
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (_GEN_373 & 3'h4 == _T_90) begin // @[InstructionMemoryCache.scala 117:47]
          buf_2_data_4 <= io_memory_response_bits_inner[63:48]; // @[InstructionMemoryCache.scala 117:47]
        end else if (_GEN_373 & 3'h4 == _T_89) begin // @[InstructionMemoryCache.scala 117:47]
          buf_2_data_4 <= io_memory_response_bits_inner[47:32]; // @[InstructionMemoryCache.scala 117:47]
        end else begin
          buf_2_data_4 <= _GEN_152;
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (_GEN_373 & 3'h5 == _T_90) begin // @[InstructionMemoryCache.scala 117:47]
          buf_2_data_5 <= io_memory_response_bits_inner[63:48]; // @[InstructionMemoryCache.scala 117:47]
        end else if (_GEN_373 & 3'h5 == _T_89) begin // @[InstructionMemoryCache.scala 117:47]
          buf_2_data_5 <= io_memory_response_bits_inner[47:32]; // @[InstructionMemoryCache.scala 117:47]
        end else begin
          buf_2_data_5 <= _GEN_153;
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (_GEN_373 & 3'h6 == _T_90) begin // @[InstructionMemoryCache.scala 117:47]
          buf_2_data_6 <= io_memory_response_bits_inner[63:48]; // @[InstructionMemoryCache.scala 117:47]
        end else if (_GEN_373 & 3'h6 == _T_89) begin // @[InstructionMemoryCache.scala 117:47]
          buf_2_data_6 <= io_memory_response_bits_inner[47:32]; // @[InstructionMemoryCache.scala 117:47]
        end else begin
          buf_2_data_6 <= _GEN_154;
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (_GEN_373 & 3'h7 == _T_90) begin // @[InstructionMemoryCache.scala 117:47]
          buf_2_data_7 <= io_memory_response_bits_inner[63:48]; // @[InstructionMemoryCache.scala 117:47]
        end else if (_GEN_373 & 3'h7 == _T_89) begin // @[InstructionMemoryCache.scala 117:47]
          buf_2_data_7 <= io_memory_response_bits_inner[47:32]; // @[InstructionMemoryCache.scala 117:47]
        end else begin
          buf_2_data_7 <= _GEN_155;
        end
      end
    end
    if (reset) begin // @[InstructionMemoryCache.scala 41:28]
      buf_3_valid <= 1'h0; // @[InstructionMemoryCache.scala 41:28]
    end else if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (readIndex) begin // @[InstructionMemoryCache.scala 121:31]
          buf_3_valid <= _GEN_231;
        end else begin
          buf_3_valid <= _GEN_99;
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (readIndex) begin // @[InstructionMemoryCache.scala 121:31]
          if (2'h3 == head) begin // @[InstructionMemoryCache.scala 124:25]
            buf_3_upper <= requested; // @[InstructionMemoryCache.scala 124:25]
          end
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (_GEN_389 & 3'h0 == _T_90) begin // @[InstructionMemoryCache.scala 117:47]
          buf_3_data_0 <= io_memory_response_bits_inner[63:48]; // @[InstructionMemoryCache.scala 117:47]
        end else if (_GEN_389 & 3'h0 == _T_89) begin // @[InstructionMemoryCache.scala 117:47]
          buf_3_data_0 <= io_memory_response_bits_inner[47:32]; // @[InstructionMemoryCache.scala 117:47]
        end else begin
          buf_3_data_0 <= _GEN_156;
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (_GEN_389 & 3'h1 == _T_90) begin // @[InstructionMemoryCache.scala 117:47]
          buf_3_data_1 <= io_memory_response_bits_inner[63:48]; // @[InstructionMemoryCache.scala 117:47]
        end else if (_GEN_389 & 3'h1 == _T_89) begin // @[InstructionMemoryCache.scala 117:47]
          buf_3_data_1 <= io_memory_response_bits_inner[47:32]; // @[InstructionMemoryCache.scala 117:47]
        end else begin
          buf_3_data_1 <= _GEN_157;
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (_GEN_389 & 3'h2 == _T_90) begin // @[InstructionMemoryCache.scala 117:47]
          buf_3_data_2 <= io_memory_response_bits_inner[63:48]; // @[InstructionMemoryCache.scala 117:47]
        end else if (_GEN_389 & 3'h2 == _T_89) begin // @[InstructionMemoryCache.scala 117:47]
          buf_3_data_2 <= io_memory_response_bits_inner[47:32]; // @[InstructionMemoryCache.scala 117:47]
        end else begin
          buf_3_data_2 <= _GEN_158;
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (_GEN_389 & 3'h3 == _T_90) begin // @[InstructionMemoryCache.scala 117:47]
          buf_3_data_3 <= io_memory_response_bits_inner[63:48]; // @[InstructionMemoryCache.scala 117:47]
        end else if (_GEN_389 & 3'h3 == _T_89) begin // @[InstructionMemoryCache.scala 117:47]
          buf_3_data_3 <= io_memory_response_bits_inner[47:32]; // @[InstructionMemoryCache.scala 117:47]
        end else begin
          buf_3_data_3 <= _GEN_159;
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (_GEN_389 & 3'h4 == _T_90) begin // @[InstructionMemoryCache.scala 117:47]
          buf_3_data_4 <= io_memory_response_bits_inner[63:48]; // @[InstructionMemoryCache.scala 117:47]
        end else if (_GEN_389 & 3'h4 == _T_89) begin // @[InstructionMemoryCache.scala 117:47]
          buf_3_data_4 <= io_memory_response_bits_inner[47:32]; // @[InstructionMemoryCache.scala 117:47]
        end else begin
          buf_3_data_4 <= _GEN_160;
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (_GEN_389 & 3'h5 == _T_90) begin // @[InstructionMemoryCache.scala 117:47]
          buf_3_data_5 <= io_memory_response_bits_inner[63:48]; // @[InstructionMemoryCache.scala 117:47]
        end else if (_GEN_389 & 3'h5 == _T_89) begin // @[InstructionMemoryCache.scala 117:47]
          buf_3_data_5 <= io_memory_response_bits_inner[47:32]; // @[InstructionMemoryCache.scala 117:47]
        end else begin
          buf_3_data_5 <= _GEN_161;
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (_GEN_389 & 3'h6 == _T_90) begin // @[InstructionMemoryCache.scala 117:47]
          buf_3_data_6 <= io_memory_response_bits_inner[63:48]; // @[InstructionMemoryCache.scala 117:47]
        end else if (_GEN_389 & 3'h6 == _T_89) begin // @[InstructionMemoryCache.scala 117:47]
          buf_3_data_6 <= io_memory_response_bits_inner[47:32]; // @[InstructionMemoryCache.scala 117:47]
        end else begin
          buf_3_data_6 <= _GEN_162;
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (_GEN_389 & 3'h7 == _T_90) begin // @[InstructionMemoryCache.scala 117:47]
          buf_3_data_7 <= io_memory_response_bits_inner[63:48]; // @[InstructionMemoryCache.scala 117:47]
        end else if (_GEN_389 & 3'h7 == _T_89) begin // @[InstructionMemoryCache.scala 117:47]
          buf_3_data_7 <= io_memory_response_bits_inner[47:32]; // @[InstructionMemoryCache.scala 117:47]
        end else begin
          buf_3_data_7 <= _GEN_163;
        end
      end
    end
    if (reset) begin // @[InstructionMemoryCache.scala 82:30]
      state <= 1'h0; // @[InstructionMemoryCache.scala 82:30]
    end else if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (readIndex) begin // @[InstructionMemoryCache.scala 121:31]
          state <= 1'h0; // @[InstructionMemoryCache.scala 122:15]
        end else begin
          state <= _GEN_75;
        end
      end else begin
        state <= _GEN_75;
      end
    end else begin
      state <= _GEN_75;
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        readIndex <= readIndex + 1'h1; // @[InstructionMemoryCache.scala 120:17]
      end else begin
        readIndex <= _GEN_77;
      end
    end else begin
      readIndex <= _GEN_77;
    end
    if (reset) begin // @[InstructionMemoryCache.scala 84:34]
      requested <= 60'h0; // @[InstructionMemoryCache.scala 84:34]
    end else if (_T_81 & ~state) begin // @[InstructionMemoryCache.scala 88:41]
      if (io_fetch_0_address_valid) begin // @[InstructionMemoryCache.scala 71:27]
        if (~_T_35) begin // @[InstructionMemoryCache.scala 72:39]
          requested <= lowerAddress[62:3]; // @[InstructionMemoryCache.scala 73:17]
        end else begin
          requested <= _GEN_72;
        end
      end else begin
        requested <= 60'h0; // @[InstructionMemoryCache.scala 43:36]
      end
    end
    if (_T_81 & ~state) begin // @[InstructionMemoryCache.scala 88:41]
      transaction_address <= tmp_transaction_address; // @[InstructionMemoryCache.scala 96:17]
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (~requestDone) begin // @[InstructionMemoryCache.scala 106:24]
        requestDone <= _GEN_86;
      end else begin
        requestDone <= _GEN_85;
      end
    end else begin
      requestDone <= _GEN_85;
    end
    if (reset) begin // @[InstructionMemoryCache.scala 104:29]
      head <= 2'h0; // @[InstructionMemoryCache.scala 104:29]
    end else if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (readIndex) begin // @[InstructionMemoryCache.scala 121:31]
          head <= _head_T_1; // @[InstructionMemoryCache.scala 125:14]
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  buf_0_valid = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  buf_0_upper = _RAND_1[59:0];
  _RAND_2 = {1{`RANDOM}};
  buf_0_data_0 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  buf_0_data_1 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  buf_0_data_2 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  buf_0_data_3 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  buf_0_data_4 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  buf_0_data_5 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  buf_0_data_6 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  buf_0_data_7 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  buf_1_valid = _RAND_10[0:0];
  _RAND_11 = {2{`RANDOM}};
  buf_1_upper = _RAND_11[59:0];
  _RAND_12 = {1{`RANDOM}};
  buf_1_data_0 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  buf_1_data_1 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  buf_1_data_2 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  buf_1_data_3 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  buf_1_data_4 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  buf_1_data_5 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  buf_1_data_6 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  buf_1_data_7 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  buf_2_valid = _RAND_20[0:0];
  _RAND_21 = {2{`RANDOM}};
  buf_2_upper = _RAND_21[59:0];
  _RAND_22 = {1{`RANDOM}};
  buf_2_data_0 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  buf_2_data_1 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  buf_2_data_2 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  buf_2_data_3 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  buf_2_data_4 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  buf_2_data_5 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  buf_2_data_6 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  buf_2_data_7 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  buf_3_valid = _RAND_30[0:0];
  _RAND_31 = {2{`RANDOM}};
  buf_3_upper = _RAND_31[59:0];
  _RAND_32 = {1{`RANDOM}};
  buf_3_data_0 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  buf_3_data_1 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  buf_3_data_2 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  buf_3_data_3 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  buf_3_data_4 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  buf_3_data_5 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  buf_3_data_6 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  buf_3_data_7 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  state = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  readIndex = _RAND_41[0:0];
  _RAND_42 = {2{`RANDOM}};
  requested = _RAND_42[59:0];
  _RAND_43 = {2{`RANDOM}};
  transaction_address = _RAND_43[63:0];
  _RAND_44 = {1{`RANDOM}};
  requestDone = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  head = _RAND_45[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module InstructionMemoryCache_1(
  input         clock,
  input         reset,
  input         io_fetch_0_address_valid,
  input  [63:0] io_fetch_0_address_bits,
  output        io_fetch_0_output_valid,
  output [31:0] io_fetch_0_output_bits,
  input         io_memory_request_ready,
  output        io_memory_request_valid,
  output [63:0] io_memory_request_bits_address,
  input         io_memory_response_valid,
  input  [63:0] io_memory_response_bits_inner
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [63:0] _RAND_42;
  reg [63:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
`endif // RANDOMIZE_REG_INIT
  reg  buf_0_valid; // @[InstructionMemoryCache.scala 41:28]
  reg [59:0] buf_0_upper; // @[InstructionMemoryCache.scala 41:28]
  reg [15:0] buf_0_data_0; // @[InstructionMemoryCache.scala 41:28]
  reg [15:0] buf_0_data_1; // @[InstructionMemoryCache.scala 41:28]
  reg [15:0] buf_0_data_2; // @[InstructionMemoryCache.scala 41:28]
  reg [15:0] buf_0_data_3; // @[InstructionMemoryCache.scala 41:28]
  reg [15:0] buf_0_data_4; // @[InstructionMemoryCache.scala 41:28]
  reg [15:0] buf_0_data_5; // @[InstructionMemoryCache.scala 41:28]
  reg [15:0] buf_0_data_6; // @[InstructionMemoryCache.scala 41:28]
  reg [15:0] buf_0_data_7; // @[InstructionMemoryCache.scala 41:28]
  reg  buf_1_valid; // @[InstructionMemoryCache.scala 41:28]
  reg [59:0] buf_1_upper; // @[InstructionMemoryCache.scala 41:28]
  reg [15:0] buf_1_data_0; // @[InstructionMemoryCache.scala 41:28]
  reg [15:0] buf_1_data_1; // @[InstructionMemoryCache.scala 41:28]
  reg [15:0] buf_1_data_2; // @[InstructionMemoryCache.scala 41:28]
  reg [15:0] buf_1_data_3; // @[InstructionMemoryCache.scala 41:28]
  reg [15:0] buf_1_data_4; // @[InstructionMemoryCache.scala 41:28]
  reg [15:0] buf_1_data_5; // @[InstructionMemoryCache.scala 41:28]
  reg [15:0] buf_1_data_6; // @[InstructionMemoryCache.scala 41:28]
  reg [15:0] buf_1_data_7; // @[InstructionMemoryCache.scala 41:28]
  reg  buf_2_valid; // @[InstructionMemoryCache.scala 41:28]
  reg [59:0] buf_2_upper; // @[InstructionMemoryCache.scala 41:28]
  reg [15:0] buf_2_data_0; // @[InstructionMemoryCache.scala 41:28]
  reg [15:0] buf_2_data_1; // @[InstructionMemoryCache.scala 41:28]
  reg [15:0] buf_2_data_2; // @[InstructionMemoryCache.scala 41:28]
  reg [15:0] buf_2_data_3; // @[InstructionMemoryCache.scala 41:28]
  reg [15:0] buf_2_data_4; // @[InstructionMemoryCache.scala 41:28]
  reg [15:0] buf_2_data_5; // @[InstructionMemoryCache.scala 41:28]
  reg [15:0] buf_2_data_6; // @[InstructionMemoryCache.scala 41:28]
  reg [15:0] buf_2_data_7; // @[InstructionMemoryCache.scala 41:28]
  reg  buf_3_valid; // @[InstructionMemoryCache.scala 41:28]
  reg [59:0] buf_3_upper; // @[InstructionMemoryCache.scala 41:28]
  reg [15:0] buf_3_data_0; // @[InstructionMemoryCache.scala 41:28]
  reg [15:0] buf_3_data_1; // @[InstructionMemoryCache.scala 41:28]
  reg [15:0] buf_3_data_2; // @[InstructionMemoryCache.scala 41:28]
  reg [15:0] buf_3_data_3; // @[InstructionMemoryCache.scala 41:28]
  reg [15:0] buf_3_data_4; // @[InstructionMemoryCache.scala 41:28]
  reg [15:0] buf_3_data_5; // @[InstructionMemoryCache.scala 41:28]
  reg [15:0] buf_3_data_6; // @[InstructionMemoryCache.scala 41:28]
  reg [15:0] buf_3_data_7; // @[InstructionMemoryCache.scala 41:28]
  wire [62:0] lowerAddress = io_fetch_0_address_bits[63:1]; // @[InstructionMemoryCache.scala 46:38]
  wire [62:0] upperAddress = lowerAddress + 63'h1; // @[InstructionMemoryCache.scala 47:37]
  wire  _T_4 = buf_0_valid & lowerAddress[62:3] == buf_0_upper; // @[InstructionMemoryCache.scala 54:34]
  wire [15:0] _GEN_1 = 3'h1 == lowerAddress[2:0] ? buf_0_data_1 : buf_0_data_0; // @[InstructionMemoryCache.scala 55:{19,19}]
  wire [15:0] _GEN_2 = 3'h2 == lowerAddress[2:0] ? buf_0_data_2 : _GEN_1; // @[InstructionMemoryCache.scala 55:{19,19}]
  wire [15:0] _GEN_3 = 3'h3 == lowerAddress[2:0] ? buf_0_data_3 : _GEN_2; // @[InstructionMemoryCache.scala 55:{19,19}]
  wire [15:0] _GEN_4 = 3'h4 == lowerAddress[2:0] ? buf_0_data_4 : _GEN_3; // @[InstructionMemoryCache.scala 55:{19,19}]
  wire [15:0] _GEN_5 = 3'h5 == lowerAddress[2:0] ? buf_0_data_5 : _GEN_4; // @[InstructionMemoryCache.scala 55:{19,19}]
  wire [15:0] _GEN_6 = 3'h6 == lowerAddress[2:0] ? buf_0_data_6 : _GEN_5; // @[InstructionMemoryCache.scala 55:{19,19}]
  wire [15:0] _GEN_7 = 3'h7 == lowerAddress[2:0] ? buf_0_data_7 : _GEN_6; // @[InstructionMemoryCache.scala 55:{19,19}]
  wire [15:0] _GEN_8 = buf_0_valid & lowerAddress[62:3] == buf_0_upper ? _GEN_7 : 16'h0; // @[InstructionMemoryCache.scala 54:70 55:19 48:32]
  wire  _T_12 = lowerAddress[62:3] == buf_1_upper; // @[InstructionMemoryCache.scala 54:57]
  wire [15:0] _GEN_10 = 3'h1 == lowerAddress[2:0] ? buf_1_data_1 : buf_1_data_0; // @[InstructionMemoryCache.scala 55:{19,19}]
  wire [15:0] _GEN_11 = 3'h2 == lowerAddress[2:0] ? buf_1_data_2 : _GEN_10; // @[InstructionMemoryCache.scala 55:{19,19}]
  wire [15:0] _GEN_12 = 3'h3 == lowerAddress[2:0] ? buf_1_data_3 : _GEN_11; // @[InstructionMemoryCache.scala 55:{19,19}]
  wire [15:0] _GEN_13 = 3'h4 == lowerAddress[2:0] ? buf_1_data_4 : _GEN_12; // @[InstructionMemoryCache.scala 55:{19,19}]
  wire [15:0] _GEN_14 = 3'h5 == lowerAddress[2:0] ? buf_1_data_5 : _GEN_13; // @[InstructionMemoryCache.scala 55:{19,19}]
  wire [15:0] _GEN_15 = 3'h6 == lowerAddress[2:0] ? buf_1_data_6 : _GEN_14; // @[InstructionMemoryCache.scala 55:{19,19}]
  wire [15:0] _GEN_16 = 3'h7 == lowerAddress[2:0] ? buf_1_data_7 : _GEN_15; // @[InstructionMemoryCache.scala 55:{19,19}]
  wire [15:0] _GEN_17 = ~(buf_0_valid & lowerAddress[62:3] == buf_0_upper) & buf_1_valid & lowerAddress[62:3] ==
    buf_1_upper ? _GEN_16 : _GEN_8; // @[InstructionMemoryCache.scala 54:70 55:19]
  wire  _T_17 = _T_4 | buf_1_valid & _T_12; // @[InstructionMemoryCache.scala 57:29]
  wire  _T_21 = lowerAddress[62:3] == buf_2_upper; // @[InstructionMemoryCache.scala 54:57]
  wire [15:0] _GEN_19 = 3'h1 == lowerAddress[2:0] ? buf_2_data_1 : buf_2_data_0; // @[InstructionMemoryCache.scala 55:{19,19}]
  wire [15:0] _GEN_20 = 3'h2 == lowerAddress[2:0] ? buf_2_data_2 : _GEN_19; // @[InstructionMemoryCache.scala 55:{19,19}]
  wire [15:0] _GEN_21 = 3'h3 == lowerAddress[2:0] ? buf_2_data_3 : _GEN_20; // @[InstructionMemoryCache.scala 55:{19,19}]
  wire [15:0] _GEN_22 = 3'h4 == lowerAddress[2:0] ? buf_2_data_4 : _GEN_21; // @[InstructionMemoryCache.scala 55:{19,19}]
  wire [15:0] _GEN_23 = 3'h5 == lowerAddress[2:0] ? buf_2_data_5 : _GEN_22; // @[InstructionMemoryCache.scala 55:{19,19}]
  wire [15:0] _GEN_24 = 3'h6 == lowerAddress[2:0] ? buf_2_data_6 : _GEN_23; // @[InstructionMemoryCache.scala 55:{19,19}]
  wire [15:0] _GEN_25 = 3'h7 == lowerAddress[2:0] ? buf_2_data_7 : _GEN_24; // @[InstructionMemoryCache.scala 55:{19,19}]
  wire [15:0] _GEN_26 = ~_T_17 & buf_2_valid & lowerAddress[62:3] == buf_2_upper ? _GEN_25 : _GEN_17; // @[InstructionMemoryCache.scala 54:70 55:19]
  wire  _T_26 = _T_4 | buf_1_valid & _T_12 | buf_2_valid & _T_21; // @[InstructionMemoryCache.scala 57:29]
  wire  _T_30 = lowerAddress[62:3] == buf_3_upper; // @[InstructionMemoryCache.scala 54:57]
  wire [15:0] _GEN_28 = 3'h1 == lowerAddress[2:0] ? buf_3_data_1 : buf_3_data_0; // @[InstructionMemoryCache.scala 55:{19,19}]
  wire [15:0] _GEN_29 = 3'h2 == lowerAddress[2:0] ? buf_3_data_2 : _GEN_28; // @[InstructionMemoryCache.scala 55:{19,19}]
  wire [15:0] _GEN_30 = 3'h3 == lowerAddress[2:0] ? buf_3_data_3 : _GEN_29; // @[InstructionMemoryCache.scala 55:{19,19}]
  wire [15:0] _GEN_31 = 3'h4 == lowerAddress[2:0] ? buf_3_data_4 : _GEN_30; // @[InstructionMemoryCache.scala 55:{19,19}]
  wire [15:0] _GEN_32 = 3'h5 == lowerAddress[2:0] ? buf_3_data_5 : _GEN_31; // @[InstructionMemoryCache.scala 55:{19,19}]
  wire [15:0] _GEN_33 = 3'h6 == lowerAddress[2:0] ? buf_3_data_6 : _GEN_32; // @[InstructionMemoryCache.scala 55:{19,19}]
  wire [15:0] _GEN_34 = 3'h7 == lowerAddress[2:0] ? buf_3_data_7 : _GEN_33; // @[InstructionMemoryCache.scala 55:{19,19}]
  wire [15:0] lowerData = ~_T_26 & buf_3_valid & lowerAddress[62:3] == buf_3_upper ? _GEN_34 : _GEN_26; // @[InstructionMemoryCache.scala 54:70 55:19]
  wire  _T_35 = _T_4 | buf_1_valid & _T_12 | buf_2_valid & _T_21 | buf_3_valid & _T_30; // @[InstructionMemoryCache.scala 57:29]
  wire  _T_40 = buf_0_valid & upperAddress[62:3] == buf_0_upper; // @[InstructionMemoryCache.scala 62:35]
  wire [15:0] _GEN_37 = 3'h1 == upperAddress[2:0] ? buf_0_data_1 : buf_0_data_0; // @[InstructionMemoryCache.scala 63:{19,19}]
  wire [15:0] _GEN_38 = 3'h2 == upperAddress[2:0] ? buf_0_data_2 : _GEN_37; // @[InstructionMemoryCache.scala 63:{19,19}]
  wire [15:0] _GEN_39 = 3'h3 == upperAddress[2:0] ? buf_0_data_3 : _GEN_38; // @[InstructionMemoryCache.scala 63:{19,19}]
  wire [15:0] _GEN_40 = 3'h4 == upperAddress[2:0] ? buf_0_data_4 : _GEN_39; // @[InstructionMemoryCache.scala 63:{19,19}]
  wire [15:0] _GEN_41 = 3'h5 == upperAddress[2:0] ? buf_0_data_5 : _GEN_40; // @[InstructionMemoryCache.scala 63:{19,19}]
  wire [15:0] _GEN_42 = 3'h6 == upperAddress[2:0] ? buf_0_data_6 : _GEN_41; // @[InstructionMemoryCache.scala 63:{19,19}]
  wire [15:0] _GEN_43 = 3'h7 == upperAddress[2:0] ? buf_0_data_7 : _GEN_42; // @[InstructionMemoryCache.scala 63:{19,19}]
  wire [15:0] _GEN_44 = buf_0_valid & upperAddress[62:3] == buf_0_upper ? _GEN_43 : 16'h0; // @[InstructionMemoryCache.scala 62:71 63:19 49:32]
  wire  _T_48 = upperAddress[62:3] == buf_1_upper; // @[InstructionMemoryCache.scala 62:58]
  wire [15:0] _GEN_46 = 3'h1 == upperAddress[2:0] ? buf_1_data_1 : buf_1_data_0; // @[InstructionMemoryCache.scala 63:{19,19}]
  wire [15:0] _GEN_47 = 3'h2 == upperAddress[2:0] ? buf_1_data_2 : _GEN_46; // @[InstructionMemoryCache.scala 63:{19,19}]
  wire [15:0] _GEN_48 = 3'h3 == upperAddress[2:0] ? buf_1_data_3 : _GEN_47; // @[InstructionMemoryCache.scala 63:{19,19}]
  wire [15:0] _GEN_49 = 3'h4 == upperAddress[2:0] ? buf_1_data_4 : _GEN_48; // @[InstructionMemoryCache.scala 63:{19,19}]
  wire [15:0] _GEN_50 = 3'h5 == upperAddress[2:0] ? buf_1_data_5 : _GEN_49; // @[InstructionMemoryCache.scala 63:{19,19}]
  wire [15:0] _GEN_51 = 3'h6 == upperAddress[2:0] ? buf_1_data_6 : _GEN_50; // @[InstructionMemoryCache.scala 63:{19,19}]
  wire [15:0] _GEN_52 = 3'h7 == upperAddress[2:0] ? buf_1_data_7 : _GEN_51; // @[InstructionMemoryCache.scala 63:{19,19}]
  wire [15:0] _GEN_53 = ~(buf_0_valid & upperAddress[62:3] == buf_0_upper) & buf_1_valid & upperAddress[62:3] ==
    buf_1_upper ? _GEN_52 : _GEN_44; // @[InstructionMemoryCache.scala 62:71 63:19]
  wire  _T_53 = _T_40 | buf_1_valid & _T_48; // @[InstructionMemoryCache.scala 65:31]
  wire  _T_57 = upperAddress[62:3] == buf_2_upper; // @[InstructionMemoryCache.scala 62:58]
  wire [15:0] _GEN_55 = 3'h1 == upperAddress[2:0] ? buf_2_data_1 : buf_2_data_0; // @[InstructionMemoryCache.scala 63:{19,19}]
  wire [15:0] _GEN_56 = 3'h2 == upperAddress[2:0] ? buf_2_data_2 : _GEN_55; // @[InstructionMemoryCache.scala 63:{19,19}]
  wire [15:0] _GEN_57 = 3'h3 == upperAddress[2:0] ? buf_2_data_3 : _GEN_56; // @[InstructionMemoryCache.scala 63:{19,19}]
  wire [15:0] _GEN_58 = 3'h4 == upperAddress[2:0] ? buf_2_data_4 : _GEN_57; // @[InstructionMemoryCache.scala 63:{19,19}]
  wire [15:0] _GEN_59 = 3'h5 == upperAddress[2:0] ? buf_2_data_5 : _GEN_58; // @[InstructionMemoryCache.scala 63:{19,19}]
  wire [15:0] _GEN_60 = 3'h6 == upperAddress[2:0] ? buf_2_data_6 : _GEN_59; // @[InstructionMemoryCache.scala 63:{19,19}]
  wire [15:0] _GEN_61 = 3'h7 == upperAddress[2:0] ? buf_2_data_7 : _GEN_60; // @[InstructionMemoryCache.scala 63:{19,19}]
  wire [15:0] _GEN_62 = ~_T_53 & buf_2_valid & upperAddress[62:3] == buf_2_upper ? _GEN_61 : _GEN_53; // @[InstructionMemoryCache.scala 62:71 63:19]
  wire  _T_62 = _T_40 | buf_1_valid & _T_48 | buf_2_valid & _T_57; // @[InstructionMemoryCache.scala 65:31]
  wire  _T_66 = upperAddress[62:3] == buf_3_upper; // @[InstructionMemoryCache.scala 62:58]
  wire [15:0] _GEN_64 = 3'h1 == upperAddress[2:0] ? buf_3_data_1 : buf_3_data_0; // @[InstructionMemoryCache.scala 63:{19,19}]
  wire [15:0] _GEN_65 = 3'h2 == upperAddress[2:0] ? buf_3_data_2 : _GEN_64; // @[InstructionMemoryCache.scala 63:{19,19}]
  wire [15:0] _GEN_66 = 3'h3 == upperAddress[2:0] ? buf_3_data_3 : _GEN_65; // @[InstructionMemoryCache.scala 63:{19,19}]
  wire [15:0] _GEN_67 = 3'h4 == upperAddress[2:0] ? buf_3_data_4 : _GEN_66; // @[InstructionMemoryCache.scala 63:{19,19}]
  wire [15:0] _GEN_68 = 3'h5 == upperAddress[2:0] ? buf_3_data_5 : _GEN_67; // @[InstructionMemoryCache.scala 63:{19,19}]
  wire [15:0] _GEN_69 = 3'h6 == upperAddress[2:0] ? buf_3_data_6 : _GEN_68; // @[InstructionMemoryCache.scala 63:{19,19}]
  wire [15:0] _GEN_70 = 3'h7 == upperAddress[2:0] ? buf_3_data_7 : _GEN_69; // @[InstructionMemoryCache.scala 63:{19,19}]
  wire [15:0] upperData = ~_T_62 & buf_3_valid & upperAddress[62:3] == buf_3_upper ? _GEN_70 : _GEN_62; // @[InstructionMemoryCache.scala 62:71 63:19]
  wire  _T_71 = _T_40 | buf_1_valid & _T_48 | buf_2_valid & _T_57 | buf_3_valid & _T_66; // @[InstructionMemoryCache.scala 65:31]
  wire  _T_72 = ~_T_35; // @[InstructionMemoryCache.scala 72:12]
  wire  _T_75 = ~_T_71; // @[InstructionMemoryCache.scala 74:18]
  wire [59:0] _GEN_72 = ~_T_71 ? upperAddress[62:3] : 60'h0; // @[InstructionMemoryCache.scala 74:46 75:17 43:36]
  wire [59:0] _GEN_73 = ~_T_35 ? lowerAddress[62:3] : _GEN_72; // @[InstructionMemoryCache.scala 72:39 73:17]
  wire [59:0] request = io_fetch_0_address_valid ? _GEN_73 : 60'h0; // @[InstructionMemoryCache.scala 71:27 43:36]
  wire  _T_81 = (_T_72 | _T_75) & io_fetch_0_address_valid; // @[InstructionMemoryCache.scala 78:60]
  reg  state; // @[InstructionMemoryCache.scala 82:30]
  reg  readIndex; // @[InstructionMemoryCache.scala 83:30]
  reg [59:0] requested; // @[InstructionMemoryCache.scala 84:34]
  reg [63:0] transaction_address; // @[InstructionMemoryCache.scala 85:32]
  reg  requestDone; // @[InstructionMemoryCache.scala 86:32]
  wire [63:0] tmp_transaction_address = {request,4'h0}; // @[Cat.scala 33:92]
  wire  _GEN_75 = _T_81 & ~state | state; // @[InstructionMemoryCache.scala 88:41 89:11 82:30]
  wire  _GEN_77 = _T_81 & ~state ? 1'h0 : readIndex; // @[InstructionMemoryCache.scala 88:41 91:15 83:30]
  wire  _GEN_85 = _T_81 & ~state ? 1'h0 : requestDone; // @[InstructionMemoryCache.scala 88:41 99:17 86:32]
  reg [1:0] head; // @[InstructionMemoryCache.scala 104:29]
  wire  _T_86 = ~requestDone; // @[InstructionMemoryCache.scala 106:10]
  wire  _GEN_86 = io_memory_request_ready | _GEN_85; // @[InstructionMemoryCache.scala 109:37 110:21]
  wire  _GEN_96 = 2'h0 == head ? 1'h0 : buf_0_valid; // @[InstructionMemoryCache.scala 115:{23,23} 41:28]
  wire  _GEN_97 = 2'h1 == head ? 1'h0 : buf_1_valid; // @[InstructionMemoryCache.scala 115:{23,23} 41:28]
  wire  _GEN_98 = 2'h2 == head ? 1'h0 : buf_2_valid; // @[InstructionMemoryCache.scala 115:{23,23} 41:28]
  wire  _GEN_99 = 2'h3 == head ? 1'h0 : buf_3_valid; // @[InstructionMemoryCache.scala 115:{23,23} 41:28]
  wire [2:0] _T_87 = {readIndex,2'h0}; // @[InstructionMemoryCache.scala 117:34]
  wire  _GEN_341 = 2'h0 == head; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [15:0] _GEN_100 = 2'h0 == head & 3'h0 == _T_87 ? io_memory_response_bits_inner[15:0] : buf_0_data_0; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [15:0] _GEN_101 = 2'h0 == head & 3'h1 == _T_87 ? io_memory_response_bits_inner[15:0] : buf_0_data_1; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [15:0] _GEN_102 = 2'h0 == head & 3'h2 == _T_87 ? io_memory_response_bits_inner[15:0] : buf_0_data_2; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [15:0] _GEN_103 = 2'h0 == head & 3'h3 == _T_87 ? io_memory_response_bits_inner[15:0] : buf_0_data_3; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [15:0] _GEN_104 = 2'h0 == head & 3'h4 == _T_87 ? io_memory_response_bits_inner[15:0] : buf_0_data_4; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [15:0] _GEN_105 = 2'h0 == head & 3'h5 == _T_87 ? io_memory_response_bits_inner[15:0] : buf_0_data_5; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [15:0] _GEN_106 = 2'h0 == head & 3'h6 == _T_87 ? io_memory_response_bits_inner[15:0] : buf_0_data_6; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [15:0] _GEN_107 = 2'h0 == head & 3'h7 == _T_87 ? io_memory_response_bits_inner[15:0] : buf_0_data_7; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire  _GEN_357 = 2'h1 == head; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [15:0] _GEN_108 = 2'h1 == head & 3'h0 == _T_87 ? io_memory_response_bits_inner[15:0] : buf_1_data_0; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [15:0] _GEN_109 = 2'h1 == head & 3'h1 == _T_87 ? io_memory_response_bits_inner[15:0] : buf_1_data_1; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [15:0] _GEN_110 = 2'h1 == head & 3'h2 == _T_87 ? io_memory_response_bits_inner[15:0] : buf_1_data_2; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [15:0] _GEN_111 = 2'h1 == head & 3'h3 == _T_87 ? io_memory_response_bits_inner[15:0] : buf_1_data_3; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [15:0] _GEN_112 = 2'h1 == head & 3'h4 == _T_87 ? io_memory_response_bits_inner[15:0] : buf_1_data_4; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [15:0] _GEN_113 = 2'h1 == head & 3'h5 == _T_87 ? io_memory_response_bits_inner[15:0] : buf_1_data_5; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [15:0] _GEN_114 = 2'h1 == head & 3'h6 == _T_87 ? io_memory_response_bits_inner[15:0] : buf_1_data_6; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [15:0] _GEN_115 = 2'h1 == head & 3'h7 == _T_87 ? io_memory_response_bits_inner[15:0] : buf_1_data_7; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire  _GEN_373 = 2'h2 == head; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [15:0] _GEN_116 = 2'h2 == head & 3'h0 == _T_87 ? io_memory_response_bits_inner[15:0] : buf_2_data_0; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [15:0] _GEN_117 = 2'h2 == head & 3'h1 == _T_87 ? io_memory_response_bits_inner[15:0] : buf_2_data_1; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [15:0] _GEN_118 = 2'h2 == head & 3'h2 == _T_87 ? io_memory_response_bits_inner[15:0] : buf_2_data_2; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [15:0] _GEN_119 = 2'h2 == head & 3'h3 == _T_87 ? io_memory_response_bits_inner[15:0] : buf_2_data_3; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [15:0] _GEN_120 = 2'h2 == head & 3'h4 == _T_87 ? io_memory_response_bits_inner[15:0] : buf_2_data_4; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [15:0] _GEN_121 = 2'h2 == head & 3'h5 == _T_87 ? io_memory_response_bits_inner[15:0] : buf_2_data_5; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [15:0] _GEN_122 = 2'h2 == head & 3'h6 == _T_87 ? io_memory_response_bits_inner[15:0] : buf_2_data_6; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [15:0] _GEN_123 = 2'h2 == head & 3'h7 == _T_87 ? io_memory_response_bits_inner[15:0] : buf_2_data_7; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire  _GEN_389 = 2'h3 == head; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [15:0] _GEN_124 = 2'h3 == head & 3'h0 == _T_87 ? io_memory_response_bits_inner[15:0] : buf_3_data_0; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [15:0] _GEN_125 = 2'h3 == head & 3'h1 == _T_87 ? io_memory_response_bits_inner[15:0] : buf_3_data_1; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [15:0] _GEN_126 = 2'h3 == head & 3'h2 == _T_87 ? io_memory_response_bits_inner[15:0] : buf_3_data_2; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [15:0] _GEN_127 = 2'h3 == head & 3'h3 == _T_87 ? io_memory_response_bits_inner[15:0] : buf_3_data_3; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [15:0] _GEN_128 = 2'h3 == head & 3'h4 == _T_87 ? io_memory_response_bits_inner[15:0] : buf_3_data_4; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [15:0] _GEN_129 = 2'h3 == head & 3'h5 == _T_87 ? io_memory_response_bits_inner[15:0] : buf_3_data_5; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [15:0] _GEN_130 = 2'h3 == head & 3'h6 == _T_87 ? io_memory_response_bits_inner[15:0] : buf_3_data_6; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [15:0] _GEN_131 = 2'h3 == head & 3'h7 == _T_87 ? io_memory_response_bits_inner[15:0] : buf_3_data_7; // @[InstructionMemoryCache.scala 117:{47,47} 41:28]
  wire [2:0] _T_88 = {readIndex,2'h1}; // @[InstructionMemoryCache.scala 117:34]
  wire [15:0] _GEN_132 = _GEN_341 & 3'h0 == _T_88 ? io_memory_response_bits_inner[31:16] : _GEN_100; // @[InstructionMemoryCache.scala 117:{47,47}]
  wire [15:0] _GEN_133 = _GEN_341 & 3'h1 == _T_88 ? io_memory_response_bits_inner[31:16] : _GEN_101; // @[InstructionMemoryCache.scala 117:{47,47}]
  wire [15:0] _GEN_134 = _GEN_341 & 3'h2 == _T_88 ? io_memory_response_bits_inner[31:16] : _GEN_102; // @[InstructionMemoryCache.scala 117:{47,47}]
  wire [15:0] _GEN_135 = _GEN_341 & 3'h3 == _T_88 ? io_memory_response_bits_inner[31:16] : _GEN_103; // @[InstructionMemoryCache.scala 117:{47,47}]
  wire [15:0] _GEN_136 = _GEN_341 & 3'h4 == _T_88 ? io_memory_response_bits_inner[31:16] : _GEN_104; // @[InstructionMemoryCache.scala 117:{47,47}]
  wire [15:0] _GEN_137 = _GEN_341 & 3'h5 == _T_88 ? io_memory_response_bits_inner[31:16] : _GEN_105; // @[InstructionMemoryCache.scala 117:{47,47}]
  wire [15:0] _GEN_138 = _GEN_341 & 3'h6 == _T_88 ? io_memory_response_bits_inner[31:16] : _GEN_106; // @[InstructionMemoryCache.scala 117:{47,47}]
  wire [15:0] _GEN_139 = _GEN_341 & 3'h7 == _T_88 ? io_memory_response_bits_inner[31:16] : _GEN_107; // @[InstructionMemoryCache.scala 117:{47,47}]
  wire [15:0] _GEN_140 = _GEN_357 & 3'h0 == _T_88 ? io_memory_response_bits_inner[31:16] : _GEN_108; // @[InstructionMemoryCache.scala 117:{47,47}]
  wire [15:0] _GEN_141 = _GEN_357 & 3'h1 == _T_88 ? io_memory_response_bits_inner[31:16] : _GEN_109; // @[InstructionMemoryCache.scala 117:{47,47}]
  wire [15:0] _GEN_142 = _GEN_357 & 3'h2 == _T_88 ? io_memory_response_bits_inner[31:16] : _GEN_110; // @[InstructionMemoryCache.scala 117:{47,47}]
  wire [15:0] _GEN_143 = _GEN_357 & 3'h3 == _T_88 ? io_memory_response_bits_inner[31:16] : _GEN_111; // @[InstructionMemoryCache.scala 117:{47,47}]
  wire [15:0] _GEN_144 = _GEN_357 & 3'h4 == _T_88 ? io_memory_response_bits_inner[31:16] : _GEN_112; // @[InstructionMemoryCache.scala 117:{47,47}]
  wire [15:0] _GEN_145 = _GEN_357 & 3'h5 == _T_88 ? io_memory_response_bits_inner[31:16] : _GEN_113; // @[InstructionMemoryCache.scala 117:{47,47}]
  wire [15:0] _GEN_146 = _GEN_357 & 3'h6 == _T_88 ? io_memory_response_bits_inner[31:16] : _GEN_114; // @[InstructionMemoryCache.scala 117:{47,47}]
  wire [15:0] _GEN_147 = _GEN_357 & 3'h7 == _T_88 ? io_memory_response_bits_inner[31:16] : _GEN_115; // @[InstructionMemoryCache.scala 117:{47,47}]
  wire [15:0] _GEN_148 = _GEN_373 & 3'h0 == _T_88 ? io_memory_response_bits_inner[31:16] : _GEN_116; // @[InstructionMemoryCache.scala 117:{47,47}]
  wire [15:0] _GEN_149 = _GEN_373 & 3'h1 == _T_88 ? io_memory_response_bits_inner[31:16] : _GEN_117; // @[InstructionMemoryCache.scala 117:{47,47}]
  wire [15:0] _GEN_150 = _GEN_373 & 3'h2 == _T_88 ? io_memory_response_bits_inner[31:16] : _GEN_118; // @[InstructionMemoryCache.scala 117:{47,47}]
  wire [15:0] _GEN_151 = _GEN_373 & 3'h3 == _T_88 ? io_memory_response_bits_inner[31:16] : _GEN_119; // @[InstructionMemoryCache.scala 117:{47,47}]
  wire [15:0] _GEN_152 = _GEN_373 & 3'h4 == _T_88 ? io_memory_response_bits_inner[31:16] : _GEN_120; // @[InstructionMemoryCache.scala 117:{47,47}]
  wire [15:0] _GEN_153 = _GEN_373 & 3'h5 == _T_88 ? io_memory_response_bits_inner[31:16] : _GEN_121; // @[InstructionMemoryCache.scala 117:{47,47}]
  wire [15:0] _GEN_154 = _GEN_373 & 3'h6 == _T_88 ? io_memory_response_bits_inner[31:16] : _GEN_122; // @[InstructionMemoryCache.scala 117:{47,47}]
  wire [15:0] _GEN_155 = _GEN_373 & 3'h7 == _T_88 ? io_memory_response_bits_inner[31:16] : _GEN_123; // @[InstructionMemoryCache.scala 117:{47,47}]
  wire [15:0] _GEN_156 = _GEN_389 & 3'h0 == _T_88 ? io_memory_response_bits_inner[31:16] : _GEN_124; // @[InstructionMemoryCache.scala 117:{47,47}]
  wire [15:0] _GEN_157 = _GEN_389 & 3'h1 == _T_88 ? io_memory_response_bits_inner[31:16] : _GEN_125; // @[InstructionMemoryCache.scala 117:{47,47}]
  wire [15:0] _GEN_158 = _GEN_389 & 3'h2 == _T_88 ? io_memory_response_bits_inner[31:16] : _GEN_126; // @[InstructionMemoryCache.scala 117:{47,47}]
  wire [15:0] _GEN_159 = _GEN_389 & 3'h3 == _T_88 ? io_memory_response_bits_inner[31:16] : _GEN_127; // @[InstructionMemoryCache.scala 117:{47,47}]
  wire [15:0] _GEN_160 = _GEN_389 & 3'h4 == _T_88 ? io_memory_response_bits_inner[31:16] : _GEN_128; // @[InstructionMemoryCache.scala 117:{47,47}]
  wire [15:0] _GEN_161 = _GEN_389 & 3'h5 == _T_88 ? io_memory_response_bits_inner[31:16] : _GEN_129; // @[InstructionMemoryCache.scala 117:{47,47}]
  wire [15:0] _GEN_162 = _GEN_389 & 3'h6 == _T_88 ? io_memory_response_bits_inner[31:16] : _GEN_130; // @[InstructionMemoryCache.scala 117:{47,47}]
  wire [15:0] _GEN_163 = _GEN_389 & 3'h7 == _T_88 ? io_memory_response_bits_inner[31:16] : _GEN_131; // @[InstructionMemoryCache.scala 117:{47,47}]
  wire [2:0] _T_89 = {readIndex,2'h2}; // @[InstructionMemoryCache.scala 117:34]
  wire [2:0] _T_90 = {readIndex,2'h3}; // @[InstructionMemoryCache.scala 117:34]
  wire  _GEN_228 = _GEN_341 | _GEN_96; // @[InstructionMemoryCache.scala 123:{25,25}]
  wire  _GEN_229 = _GEN_357 | _GEN_97; // @[InstructionMemoryCache.scala 123:{25,25}]
  wire  _GEN_230 = _GEN_373 | _GEN_98; // @[InstructionMemoryCache.scala 123:{25,25}]
  wire  _GEN_231 = _GEN_389 | _GEN_99; // @[InstructionMemoryCache.scala 123:{25,25}]
  wire [1:0] _head_T_1 = head + 2'h1; // @[InstructionMemoryCache.scala 125:22]
  assign io_fetch_0_output_valid = _T_35 & _T_71; // @[InstructionMemoryCache.scala 68:33]
  assign io_fetch_0_output_bits = {upperData,lowerData}; // @[InstructionMemoryCache.scala 69:32]
  assign io_memory_request_valid = state & _T_86; // @[InstructionMemoryCache.scala 102:27 105:30]
  assign io_memory_request_bits_address = transaction_address; // @[InstructionMemoryCache.scala 106:24 108:30]
  always @(posedge clock) begin
    if (reset) begin // @[InstructionMemoryCache.scala 41:28]
      buf_0_valid <= 1'h0; // @[InstructionMemoryCache.scala 41:28]
    end else if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (readIndex) begin // @[InstructionMemoryCache.scala 121:31]
          buf_0_valid <= _GEN_228;
        end else begin
          buf_0_valid <= _GEN_96;
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (readIndex) begin // @[InstructionMemoryCache.scala 121:31]
          if (2'h0 == head) begin // @[InstructionMemoryCache.scala 124:25]
            buf_0_upper <= requested; // @[InstructionMemoryCache.scala 124:25]
          end
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (_GEN_341 & 3'h0 == _T_90) begin // @[InstructionMemoryCache.scala 117:47]
          buf_0_data_0 <= io_memory_response_bits_inner[63:48]; // @[InstructionMemoryCache.scala 117:47]
        end else if (_GEN_341 & 3'h0 == _T_89) begin // @[InstructionMemoryCache.scala 117:47]
          buf_0_data_0 <= io_memory_response_bits_inner[47:32]; // @[InstructionMemoryCache.scala 117:47]
        end else begin
          buf_0_data_0 <= _GEN_132;
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (_GEN_341 & 3'h1 == _T_90) begin // @[InstructionMemoryCache.scala 117:47]
          buf_0_data_1 <= io_memory_response_bits_inner[63:48]; // @[InstructionMemoryCache.scala 117:47]
        end else if (_GEN_341 & 3'h1 == _T_89) begin // @[InstructionMemoryCache.scala 117:47]
          buf_0_data_1 <= io_memory_response_bits_inner[47:32]; // @[InstructionMemoryCache.scala 117:47]
        end else begin
          buf_0_data_1 <= _GEN_133;
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (_GEN_341 & 3'h2 == _T_90) begin // @[InstructionMemoryCache.scala 117:47]
          buf_0_data_2 <= io_memory_response_bits_inner[63:48]; // @[InstructionMemoryCache.scala 117:47]
        end else if (_GEN_341 & 3'h2 == _T_89) begin // @[InstructionMemoryCache.scala 117:47]
          buf_0_data_2 <= io_memory_response_bits_inner[47:32]; // @[InstructionMemoryCache.scala 117:47]
        end else begin
          buf_0_data_2 <= _GEN_134;
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (_GEN_341 & 3'h3 == _T_90) begin // @[InstructionMemoryCache.scala 117:47]
          buf_0_data_3 <= io_memory_response_bits_inner[63:48]; // @[InstructionMemoryCache.scala 117:47]
        end else if (_GEN_341 & 3'h3 == _T_89) begin // @[InstructionMemoryCache.scala 117:47]
          buf_0_data_3 <= io_memory_response_bits_inner[47:32]; // @[InstructionMemoryCache.scala 117:47]
        end else begin
          buf_0_data_3 <= _GEN_135;
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (_GEN_341 & 3'h4 == _T_90) begin // @[InstructionMemoryCache.scala 117:47]
          buf_0_data_4 <= io_memory_response_bits_inner[63:48]; // @[InstructionMemoryCache.scala 117:47]
        end else if (_GEN_341 & 3'h4 == _T_89) begin // @[InstructionMemoryCache.scala 117:47]
          buf_0_data_4 <= io_memory_response_bits_inner[47:32]; // @[InstructionMemoryCache.scala 117:47]
        end else begin
          buf_0_data_4 <= _GEN_136;
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (_GEN_341 & 3'h5 == _T_90) begin // @[InstructionMemoryCache.scala 117:47]
          buf_0_data_5 <= io_memory_response_bits_inner[63:48]; // @[InstructionMemoryCache.scala 117:47]
        end else if (_GEN_341 & 3'h5 == _T_89) begin // @[InstructionMemoryCache.scala 117:47]
          buf_0_data_5 <= io_memory_response_bits_inner[47:32]; // @[InstructionMemoryCache.scala 117:47]
        end else begin
          buf_0_data_5 <= _GEN_137;
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (_GEN_341 & 3'h6 == _T_90) begin // @[InstructionMemoryCache.scala 117:47]
          buf_0_data_6 <= io_memory_response_bits_inner[63:48]; // @[InstructionMemoryCache.scala 117:47]
        end else if (_GEN_341 & 3'h6 == _T_89) begin // @[InstructionMemoryCache.scala 117:47]
          buf_0_data_6 <= io_memory_response_bits_inner[47:32]; // @[InstructionMemoryCache.scala 117:47]
        end else begin
          buf_0_data_6 <= _GEN_138;
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (_GEN_341 & 3'h7 == _T_90) begin // @[InstructionMemoryCache.scala 117:47]
          buf_0_data_7 <= io_memory_response_bits_inner[63:48]; // @[InstructionMemoryCache.scala 117:47]
        end else if (_GEN_341 & 3'h7 == _T_89) begin // @[InstructionMemoryCache.scala 117:47]
          buf_0_data_7 <= io_memory_response_bits_inner[47:32]; // @[InstructionMemoryCache.scala 117:47]
        end else begin
          buf_0_data_7 <= _GEN_139;
        end
      end
    end
    if (reset) begin // @[InstructionMemoryCache.scala 41:28]
      buf_1_valid <= 1'h0; // @[InstructionMemoryCache.scala 41:28]
    end else if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (readIndex) begin // @[InstructionMemoryCache.scala 121:31]
          buf_1_valid <= _GEN_229;
        end else begin
          buf_1_valid <= _GEN_97;
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (readIndex) begin // @[InstructionMemoryCache.scala 121:31]
          if (2'h1 == head) begin // @[InstructionMemoryCache.scala 124:25]
            buf_1_upper <= requested; // @[InstructionMemoryCache.scala 124:25]
          end
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (_GEN_357 & 3'h0 == _T_90) begin // @[InstructionMemoryCache.scala 117:47]
          buf_1_data_0 <= io_memory_response_bits_inner[63:48]; // @[InstructionMemoryCache.scala 117:47]
        end else if (_GEN_357 & 3'h0 == _T_89) begin // @[InstructionMemoryCache.scala 117:47]
          buf_1_data_0 <= io_memory_response_bits_inner[47:32]; // @[InstructionMemoryCache.scala 117:47]
        end else begin
          buf_1_data_0 <= _GEN_140;
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (_GEN_357 & 3'h1 == _T_90) begin // @[InstructionMemoryCache.scala 117:47]
          buf_1_data_1 <= io_memory_response_bits_inner[63:48]; // @[InstructionMemoryCache.scala 117:47]
        end else if (_GEN_357 & 3'h1 == _T_89) begin // @[InstructionMemoryCache.scala 117:47]
          buf_1_data_1 <= io_memory_response_bits_inner[47:32]; // @[InstructionMemoryCache.scala 117:47]
        end else begin
          buf_1_data_1 <= _GEN_141;
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (_GEN_357 & 3'h2 == _T_90) begin // @[InstructionMemoryCache.scala 117:47]
          buf_1_data_2 <= io_memory_response_bits_inner[63:48]; // @[InstructionMemoryCache.scala 117:47]
        end else if (_GEN_357 & 3'h2 == _T_89) begin // @[InstructionMemoryCache.scala 117:47]
          buf_1_data_2 <= io_memory_response_bits_inner[47:32]; // @[InstructionMemoryCache.scala 117:47]
        end else begin
          buf_1_data_2 <= _GEN_142;
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (_GEN_357 & 3'h3 == _T_90) begin // @[InstructionMemoryCache.scala 117:47]
          buf_1_data_3 <= io_memory_response_bits_inner[63:48]; // @[InstructionMemoryCache.scala 117:47]
        end else if (_GEN_357 & 3'h3 == _T_89) begin // @[InstructionMemoryCache.scala 117:47]
          buf_1_data_3 <= io_memory_response_bits_inner[47:32]; // @[InstructionMemoryCache.scala 117:47]
        end else begin
          buf_1_data_3 <= _GEN_143;
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (_GEN_357 & 3'h4 == _T_90) begin // @[InstructionMemoryCache.scala 117:47]
          buf_1_data_4 <= io_memory_response_bits_inner[63:48]; // @[InstructionMemoryCache.scala 117:47]
        end else if (_GEN_357 & 3'h4 == _T_89) begin // @[InstructionMemoryCache.scala 117:47]
          buf_1_data_4 <= io_memory_response_bits_inner[47:32]; // @[InstructionMemoryCache.scala 117:47]
        end else begin
          buf_1_data_4 <= _GEN_144;
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (_GEN_357 & 3'h5 == _T_90) begin // @[InstructionMemoryCache.scala 117:47]
          buf_1_data_5 <= io_memory_response_bits_inner[63:48]; // @[InstructionMemoryCache.scala 117:47]
        end else if (_GEN_357 & 3'h5 == _T_89) begin // @[InstructionMemoryCache.scala 117:47]
          buf_1_data_5 <= io_memory_response_bits_inner[47:32]; // @[InstructionMemoryCache.scala 117:47]
        end else begin
          buf_1_data_5 <= _GEN_145;
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (_GEN_357 & 3'h6 == _T_90) begin // @[InstructionMemoryCache.scala 117:47]
          buf_1_data_6 <= io_memory_response_bits_inner[63:48]; // @[InstructionMemoryCache.scala 117:47]
        end else if (_GEN_357 & 3'h6 == _T_89) begin // @[InstructionMemoryCache.scala 117:47]
          buf_1_data_6 <= io_memory_response_bits_inner[47:32]; // @[InstructionMemoryCache.scala 117:47]
        end else begin
          buf_1_data_6 <= _GEN_146;
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (_GEN_357 & 3'h7 == _T_90) begin // @[InstructionMemoryCache.scala 117:47]
          buf_1_data_7 <= io_memory_response_bits_inner[63:48]; // @[InstructionMemoryCache.scala 117:47]
        end else if (_GEN_357 & 3'h7 == _T_89) begin // @[InstructionMemoryCache.scala 117:47]
          buf_1_data_7 <= io_memory_response_bits_inner[47:32]; // @[InstructionMemoryCache.scala 117:47]
        end else begin
          buf_1_data_7 <= _GEN_147;
        end
      end
    end
    if (reset) begin // @[InstructionMemoryCache.scala 41:28]
      buf_2_valid <= 1'h0; // @[InstructionMemoryCache.scala 41:28]
    end else if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (readIndex) begin // @[InstructionMemoryCache.scala 121:31]
          buf_2_valid <= _GEN_230;
        end else begin
          buf_2_valid <= _GEN_98;
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (readIndex) begin // @[InstructionMemoryCache.scala 121:31]
          if (2'h2 == head) begin // @[InstructionMemoryCache.scala 124:25]
            buf_2_upper <= requested; // @[InstructionMemoryCache.scala 124:25]
          end
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (_GEN_373 & 3'h0 == _T_90) begin // @[InstructionMemoryCache.scala 117:47]
          buf_2_data_0 <= io_memory_response_bits_inner[63:48]; // @[InstructionMemoryCache.scala 117:47]
        end else if (_GEN_373 & 3'h0 == _T_89) begin // @[InstructionMemoryCache.scala 117:47]
          buf_2_data_0 <= io_memory_response_bits_inner[47:32]; // @[InstructionMemoryCache.scala 117:47]
        end else begin
          buf_2_data_0 <= _GEN_148;
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (_GEN_373 & 3'h1 == _T_90) begin // @[InstructionMemoryCache.scala 117:47]
          buf_2_data_1 <= io_memory_response_bits_inner[63:48]; // @[InstructionMemoryCache.scala 117:47]
        end else if (_GEN_373 & 3'h1 == _T_89) begin // @[InstructionMemoryCache.scala 117:47]
          buf_2_data_1 <= io_memory_response_bits_inner[47:32]; // @[InstructionMemoryCache.scala 117:47]
        end else begin
          buf_2_data_1 <= _GEN_149;
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (_GEN_373 & 3'h2 == _T_90) begin // @[InstructionMemoryCache.scala 117:47]
          buf_2_data_2 <= io_memory_response_bits_inner[63:48]; // @[InstructionMemoryCache.scala 117:47]
        end else if (_GEN_373 & 3'h2 == _T_89) begin // @[InstructionMemoryCache.scala 117:47]
          buf_2_data_2 <= io_memory_response_bits_inner[47:32]; // @[InstructionMemoryCache.scala 117:47]
        end else begin
          buf_2_data_2 <= _GEN_150;
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (_GEN_373 & 3'h3 == _T_90) begin // @[InstructionMemoryCache.scala 117:47]
          buf_2_data_3 <= io_memory_response_bits_inner[63:48]; // @[InstructionMemoryCache.scala 117:47]
        end else if (_GEN_373 & 3'h3 == _T_89) begin // @[InstructionMemoryCache.scala 117:47]
          buf_2_data_3 <= io_memory_response_bits_inner[47:32]; // @[InstructionMemoryCache.scala 117:47]
        end else begin
          buf_2_data_3 <= _GEN_151;
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (_GEN_373 & 3'h4 == _T_90) begin // @[InstructionMemoryCache.scala 117:47]
          buf_2_data_4 <= io_memory_response_bits_inner[63:48]; // @[InstructionMemoryCache.scala 117:47]
        end else if (_GEN_373 & 3'h4 == _T_89) begin // @[InstructionMemoryCache.scala 117:47]
          buf_2_data_4 <= io_memory_response_bits_inner[47:32]; // @[InstructionMemoryCache.scala 117:47]
        end else begin
          buf_2_data_4 <= _GEN_152;
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (_GEN_373 & 3'h5 == _T_90) begin // @[InstructionMemoryCache.scala 117:47]
          buf_2_data_5 <= io_memory_response_bits_inner[63:48]; // @[InstructionMemoryCache.scala 117:47]
        end else if (_GEN_373 & 3'h5 == _T_89) begin // @[InstructionMemoryCache.scala 117:47]
          buf_2_data_5 <= io_memory_response_bits_inner[47:32]; // @[InstructionMemoryCache.scala 117:47]
        end else begin
          buf_2_data_5 <= _GEN_153;
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (_GEN_373 & 3'h6 == _T_90) begin // @[InstructionMemoryCache.scala 117:47]
          buf_2_data_6 <= io_memory_response_bits_inner[63:48]; // @[InstructionMemoryCache.scala 117:47]
        end else if (_GEN_373 & 3'h6 == _T_89) begin // @[InstructionMemoryCache.scala 117:47]
          buf_2_data_6 <= io_memory_response_bits_inner[47:32]; // @[InstructionMemoryCache.scala 117:47]
        end else begin
          buf_2_data_6 <= _GEN_154;
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (_GEN_373 & 3'h7 == _T_90) begin // @[InstructionMemoryCache.scala 117:47]
          buf_2_data_7 <= io_memory_response_bits_inner[63:48]; // @[InstructionMemoryCache.scala 117:47]
        end else if (_GEN_373 & 3'h7 == _T_89) begin // @[InstructionMemoryCache.scala 117:47]
          buf_2_data_7 <= io_memory_response_bits_inner[47:32]; // @[InstructionMemoryCache.scala 117:47]
        end else begin
          buf_2_data_7 <= _GEN_155;
        end
      end
    end
    if (reset) begin // @[InstructionMemoryCache.scala 41:28]
      buf_3_valid <= 1'h0; // @[InstructionMemoryCache.scala 41:28]
    end else if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (readIndex) begin // @[InstructionMemoryCache.scala 121:31]
          buf_3_valid <= _GEN_231;
        end else begin
          buf_3_valid <= _GEN_99;
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (readIndex) begin // @[InstructionMemoryCache.scala 121:31]
          if (2'h3 == head) begin // @[InstructionMemoryCache.scala 124:25]
            buf_3_upper <= requested; // @[InstructionMemoryCache.scala 124:25]
          end
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (_GEN_389 & 3'h0 == _T_90) begin // @[InstructionMemoryCache.scala 117:47]
          buf_3_data_0 <= io_memory_response_bits_inner[63:48]; // @[InstructionMemoryCache.scala 117:47]
        end else if (_GEN_389 & 3'h0 == _T_89) begin // @[InstructionMemoryCache.scala 117:47]
          buf_3_data_0 <= io_memory_response_bits_inner[47:32]; // @[InstructionMemoryCache.scala 117:47]
        end else begin
          buf_3_data_0 <= _GEN_156;
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (_GEN_389 & 3'h1 == _T_90) begin // @[InstructionMemoryCache.scala 117:47]
          buf_3_data_1 <= io_memory_response_bits_inner[63:48]; // @[InstructionMemoryCache.scala 117:47]
        end else if (_GEN_389 & 3'h1 == _T_89) begin // @[InstructionMemoryCache.scala 117:47]
          buf_3_data_1 <= io_memory_response_bits_inner[47:32]; // @[InstructionMemoryCache.scala 117:47]
        end else begin
          buf_3_data_1 <= _GEN_157;
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (_GEN_389 & 3'h2 == _T_90) begin // @[InstructionMemoryCache.scala 117:47]
          buf_3_data_2 <= io_memory_response_bits_inner[63:48]; // @[InstructionMemoryCache.scala 117:47]
        end else if (_GEN_389 & 3'h2 == _T_89) begin // @[InstructionMemoryCache.scala 117:47]
          buf_3_data_2 <= io_memory_response_bits_inner[47:32]; // @[InstructionMemoryCache.scala 117:47]
        end else begin
          buf_3_data_2 <= _GEN_158;
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (_GEN_389 & 3'h3 == _T_90) begin // @[InstructionMemoryCache.scala 117:47]
          buf_3_data_3 <= io_memory_response_bits_inner[63:48]; // @[InstructionMemoryCache.scala 117:47]
        end else if (_GEN_389 & 3'h3 == _T_89) begin // @[InstructionMemoryCache.scala 117:47]
          buf_3_data_3 <= io_memory_response_bits_inner[47:32]; // @[InstructionMemoryCache.scala 117:47]
        end else begin
          buf_3_data_3 <= _GEN_159;
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (_GEN_389 & 3'h4 == _T_90) begin // @[InstructionMemoryCache.scala 117:47]
          buf_3_data_4 <= io_memory_response_bits_inner[63:48]; // @[InstructionMemoryCache.scala 117:47]
        end else if (_GEN_389 & 3'h4 == _T_89) begin // @[InstructionMemoryCache.scala 117:47]
          buf_3_data_4 <= io_memory_response_bits_inner[47:32]; // @[InstructionMemoryCache.scala 117:47]
        end else begin
          buf_3_data_4 <= _GEN_160;
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (_GEN_389 & 3'h5 == _T_90) begin // @[InstructionMemoryCache.scala 117:47]
          buf_3_data_5 <= io_memory_response_bits_inner[63:48]; // @[InstructionMemoryCache.scala 117:47]
        end else if (_GEN_389 & 3'h5 == _T_89) begin // @[InstructionMemoryCache.scala 117:47]
          buf_3_data_5 <= io_memory_response_bits_inner[47:32]; // @[InstructionMemoryCache.scala 117:47]
        end else begin
          buf_3_data_5 <= _GEN_161;
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (_GEN_389 & 3'h6 == _T_90) begin // @[InstructionMemoryCache.scala 117:47]
          buf_3_data_6 <= io_memory_response_bits_inner[63:48]; // @[InstructionMemoryCache.scala 117:47]
        end else if (_GEN_389 & 3'h6 == _T_89) begin // @[InstructionMemoryCache.scala 117:47]
          buf_3_data_6 <= io_memory_response_bits_inner[47:32]; // @[InstructionMemoryCache.scala 117:47]
        end else begin
          buf_3_data_6 <= _GEN_162;
        end
      end
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (_GEN_389 & 3'h7 == _T_90) begin // @[InstructionMemoryCache.scala 117:47]
          buf_3_data_7 <= io_memory_response_bits_inner[63:48]; // @[InstructionMemoryCache.scala 117:47]
        end else if (_GEN_389 & 3'h7 == _T_89) begin // @[InstructionMemoryCache.scala 117:47]
          buf_3_data_7 <= io_memory_response_bits_inner[47:32]; // @[InstructionMemoryCache.scala 117:47]
        end else begin
          buf_3_data_7 <= _GEN_163;
        end
      end
    end
    if (reset) begin // @[InstructionMemoryCache.scala 82:30]
      state <= 1'h0; // @[InstructionMemoryCache.scala 82:30]
    end else if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (readIndex) begin // @[InstructionMemoryCache.scala 121:31]
          state <= 1'h0; // @[InstructionMemoryCache.scala 122:15]
        end else begin
          state <= _GEN_75;
        end
      end else begin
        state <= _GEN_75;
      end
    end else begin
      state <= _GEN_75;
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        readIndex <= readIndex + 1'h1; // @[InstructionMemoryCache.scala 120:17]
      end else begin
        readIndex <= _GEN_77;
      end
    end else begin
      readIndex <= _GEN_77;
    end
    if (reset) begin // @[InstructionMemoryCache.scala 84:34]
      requested <= 60'h0; // @[InstructionMemoryCache.scala 84:34]
    end else if (_T_81 & ~state) begin // @[InstructionMemoryCache.scala 88:41]
      if (io_fetch_0_address_valid) begin // @[InstructionMemoryCache.scala 71:27]
        if (~_T_35) begin // @[InstructionMemoryCache.scala 72:39]
          requested <= lowerAddress[62:3]; // @[InstructionMemoryCache.scala 73:17]
        end else begin
          requested <= _GEN_72;
        end
      end else begin
        requested <= 60'h0; // @[InstructionMemoryCache.scala 43:36]
      end
    end
    if (_T_81 & ~state) begin // @[InstructionMemoryCache.scala 88:41]
      transaction_address <= tmp_transaction_address; // @[InstructionMemoryCache.scala 96:17]
    end
    if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (~requestDone) begin // @[InstructionMemoryCache.scala 106:24]
        requestDone <= _GEN_86;
      end else begin
        requestDone <= _GEN_85;
      end
    end else begin
      requestDone <= _GEN_85;
    end
    if (reset) begin // @[InstructionMemoryCache.scala 104:29]
      head <= 2'h0; // @[InstructionMemoryCache.scala 104:29]
    end else if (state) begin // @[InstructionMemoryCache.scala 105:30]
      if (io_memory_response_valid) begin // @[InstructionMemoryCache.scala 114:36]
        if (readIndex) begin // @[InstructionMemoryCache.scala 121:31]
          head <= _head_T_1; // @[InstructionMemoryCache.scala 125:14]
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  buf_0_valid = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  buf_0_upper = _RAND_1[59:0];
  _RAND_2 = {1{`RANDOM}};
  buf_0_data_0 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  buf_0_data_1 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  buf_0_data_2 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  buf_0_data_3 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  buf_0_data_4 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  buf_0_data_5 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  buf_0_data_6 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  buf_0_data_7 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  buf_1_valid = _RAND_10[0:0];
  _RAND_11 = {2{`RANDOM}};
  buf_1_upper = _RAND_11[59:0];
  _RAND_12 = {1{`RANDOM}};
  buf_1_data_0 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  buf_1_data_1 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  buf_1_data_2 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  buf_1_data_3 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  buf_1_data_4 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  buf_1_data_5 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  buf_1_data_6 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  buf_1_data_7 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  buf_2_valid = _RAND_20[0:0];
  _RAND_21 = {2{`RANDOM}};
  buf_2_upper = _RAND_21[59:0];
  _RAND_22 = {1{`RANDOM}};
  buf_2_data_0 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  buf_2_data_1 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  buf_2_data_2 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  buf_2_data_3 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  buf_2_data_4 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  buf_2_data_5 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  buf_2_data_6 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  buf_2_data_7 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  buf_3_valid = _RAND_30[0:0];
  _RAND_31 = {2{`RANDOM}};
  buf_3_upper = _RAND_31[59:0];
  _RAND_32 = {1{`RANDOM}};
  buf_3_data_0 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  buf_3_data_1 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  buf_3_data_2 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  buf_3_data_3 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  buf_3_data_4 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  buf_3_data_5 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  buf_3_data_6 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  buf_3_data_7 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  state = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  readIndex = _RAND_41[0:0];
  _RAND_42 = {2{`RANDOM}};
  requested = _RAND_42[59:0];
  _RAND_43 = {2{`RANDOM}};
  transaction_address = _RAND_43[63:0];
  _RAND_44 = {1{`RANDOM}};
  requestDone = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  head = _RAND_45[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CheckBranch(
  input  [31:0] io_instruction,
  output [3:0]  io_branchType,
  output [20:0] io_offset
);
  wire [6:0] opcode = io_instruction[6:0]; // @[CheckBranch.scala 22:30]
  wire [2:0] funct3 = io_instruction[14:12]; // @[CheckBranch.scala 25:30]
  wire [2:0] _io_offset_T_2 = io_instruction[15:13] & 3'h3; // @[CheckBranch.scala 34:32]
  wire  _io_offset_T_3 = 3'h1 == _io_offset_T_2; // @[CheckBranch.scala 34:32]
  wire [11:0] _io_offset_T_13 = {io_instruction[12],io_instruction[8],io_instruction[10:9],io_instruction[6],
    io_instruction[7],io_instruction[2],io_instruction[11],io_instruction[5:3],1'h0}; // @[CheckBranch.scala 45:11]
  wire [11:0] _io_offset_T_14 = _io_offset_T_3 ? $signed(_io_offset_T_13) : $signed(12'sh2); // @[CheckBranch.scala 33:21]
  wire  _io_offset_T_18 = io_instruction[11:7] != 5'h0; // @[CheckBranch.scala 52:35]
  wire  _io_offset_T_19 = io_instruction[15:13] == 3'h4 & _io_offset_T_18; // @[CheckBranch.scala 51:48]
  wire  _io_offset_T_21 = io_instruction[6:2] == 5'h0; // @[CheckBranch.scala 53:34]
  wire  _io_offset_T_22 = _io_offset_T_19 & _io_offset_T_21; // @[CheckBranch.scala 52:43]
  wire  _io_offset_T_26 = io_instruction[11:7] == 5'h0; // @[CheckBranch.scala 55:35]
  wire  _io_offset_T_27 = io_instruction[15:12] == 4'h9 & _io_offset_T_26; // @[CheckBranch.scala 54:49]
  wire  _io_offset_T_30 = _io_offset_T_27 & _io_offset_T_21; // @[CheckBranch.scala 55:43]
  wire [2:0] _io_offset_T_31 = _io_offset_T_30 ? $signed(3'sh0) : $signed(3'sh2); // @[Mux.scala 101:16]
  wire [2:0] _io_offset_T_32 = _io_offset_T_22 ? $signed(3'sh0) : $signed(_io_offset_T_31); // @[Mux.scala 101:16]
  wire [12:0] _io_offset_T_35 = {io_instruction[31:20],1'h0}; // @[CheckBranch.scala 64:65]
  wire [20:0] _io_offset_T_41 = {io_instruction[31],io_instruction[19:12],io_instruction[20],io_instruction[30:21],1'h0}
    ; // @[CheckBranch.scala 72:13]
  wire [12:0] _io_offset_T_43 = 7'h67 == opcode ? $signed(_io_offset_T_35) : $signed(13'sh4); // @[Mux.scala 81:58]
  wire [20:0] _io_offset_T_45 = 7'h6f == opcode ? $signed(_io_offset_T_41) : $signed({{8{_io_offset_T_43[12]}},
    _io_offset_T_43}); // @[Mux.scala 81:58]
  wire [20:0] _io_offset_T_47 = 7'h63 == opcode ? $signed(21'sh4) : $signed(_io_offset_T_45); // @[Mux.scala 81:58]
  wire [20:0] _io_offset_T_49 = 7'hf == opcode ? $signed(21'sh4) : $signed(_io_offset_T_47); // @[Mux.scala 81:58]
  wire [11:0] _io_offset_T_51 = 2'h1 == opcode[1:0] ? $signed(_io_offset_T_14) : $signed(12'sh2); // @[Mux.scala 81:58]
  wire [11:0] _io_offset_T_53 = 2'h2 == opcode[1:0] ? $signed({{9{_io_offset_T_32[2]}},_io_offset_T_32}) : $signed(
    _io_offset_T_51); // @[Mux.scala 81:58]
  wire  _io_branchType_T_3 = 3'h5 == io_instruction[15:13]; // @[CheckBranch.scala 91:35]
  wire [2:0] _io_branchType_T_5 = io_instruction[15:13] & 3'h6; // @[CheckBranch.scala 92:35]
  wire  _io_branchType_T_6 = 3'h6 == _io_branchType_T_5; // @[CheckBranch.scala 92:35]
  wire [1:0] _io_branchType_T_7 = _io_branchType_T_6 ? 2'h2 : 2'h1; // @[Mux.scala 101:16]
  wire [1:0] _io_branchType_T_8 = _io_branchType_T_3 ? 2'h3 : _io_branchType_T_7; // @[Mux.scala 101:16]
  wire [3:0] _io_branchType_T_25 = _io_offset_T_30 ? 4'h8 : 4'h1; // @[Mux.scala 101:16]
  wire [3:0] _io_branchType_T_26 = _io_offset_T_22 ? 4'h4 : _io_branchType_T_25; // @[Mux.scala 101:16]
  wire [2:0] _io_branchType_T_28 = io_instruction[12] ? 3'h6 : 3'h5; // @[CheckBranch.scala 117:30]
  wire [2:0] _io_branchType_T_30 = funct3 == 3'h0 ? 3'h7 : 3'h0; // @[CheckBranch.scala 122:30]
  wire [2:0] _io_branchType_T_32 = 7'h67 == opcode ? 3'h4 : 3'h0; // @[Mux.scala 81:58]
  wire [2:0] _io_branchType_T_34 = 7'h6f == opcode ? 3'h3 : _io_branchType_T_32; // @[Mux.scala 81:58]
  wire [2:0] _io_branchType_T_36 = 7'h63 == opcode ? 3'h2 : _io_branchType_T_34; // @[Mux.scala 81:58]
  wire [2:0] _io_branchType_T_38 = 7'hf == opcode ? _io_branchType_T_28 : _io_branchType_T_36; // @[Mux.scala 81:58]
  wire [2:0] _io_branchType_T_40 = 7'h73 == opcode ? _io_branchType_T_30 : _io_branchType_T_38; // @[Mux.scala 81:58]
  wire [1:0] _io_branchType_T_42 = 2'h1 == opcode[1:0] ? _io_branchType_T_8 : 2'h1; // @[Mux.scala 81:58]
  wire [3:0] _io_branchType_T_44 = 2'h2 == opcode[1:0] ? _io_branchType_T_26 : {{2'd0}, _io_branchType_T_42}; // @[Mux.scala 81:58]
  assign io_branchType = 2'h3 == opcode[1:0] ? {{1'd0}, _io_branchType_T_40} : _io_branchType_T_44; // @[Mux.scala 81:58]
  assign io_offset = 2'h3 == opcode[1:0] ? $signed(_io_offset_T_49) : $signed({{9{_io_offset_T_53[11]}},_io_offset_T_53}
    ); // @[Mux.scala 81:58]
endmodule
module Fetch(
  input         clock,
  input         reset,
  output        io_cache_0_address_valid,
  output [63:0] io_cache_0_address_bits,
  input         io_cache_0_output_valid,
  input  [31:0] io_cache_0_output_bits,
  input         io_reorderBufferEmpty,
  input         io_loadStoreQueueEmpty,
  input         io_collectedBranchAddresses_addresses_valid,
  input         io_collectedBranchAddresses_addresses_bits_threadId,
  input  [63:0] io_collectedBranchAddresses_addresses_bits_programCounterOffset,
  input         io_fetchBuffer_toBuffer_0_ready,
  output        io_fetchBuffer_toBuffer_0_valid,
  output [31:0] io_fetchBuffer_toBuffer_0_bits_instruction,
  output [63:0] io_fetchBuffer_toBuffer_0_bits_programCounter,
  input         io_fetchBuffer_empty,
  input  [63:0] io_csr_mtvec,
  input  [63:0] io_csr_mepc,
  input  [63:0] io_csr_mcause,
  input         io_csrReservationStationEmpty,
  input         io_isError
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] checkBranches_0_io_instruction; // @[Fetch.scala 54:63]
  wire [3:0] checkBranches_0_io_branchType; // @[Fetch.scala 54:63]
  wire [20:0] checkBranches_0_io_offset; // @[Fetch.scala 54:63]
  reg [63:0] pc; // @[Fetch.scala 57:19]
  reg [2:0] waiting; // @[Fetch.scala 60:24]
  wire  instructionValid = io_cache_0_output_valid & waiting == 3'h0; // @[Fetch.scala 76:47]
  wire  _T = waiting != 3'h0; // @[Fetch.scala 85:16]
  wire  _T_1 = ~io_fetchBuffer_toBuffer_0_ready; // @[Fetch.scala 85:42]
  wire  _T_4 = waiting != 3'h0 | ~io_fetchBuffer_toBuffer_0_ready | ~instructionValid; // @[Fetch.scala 85:57]
  wire [3:0] _T_5 = checkBranches_0_io_branchType; // @[Fetch.scala 88:30]
  wire  _T_11 = $signed(checkBranches_0_io_offset) == 21'sh0; // @[Fetch.scala 96:30]
  wire [2:0] _T_12 = _T_11 ? 3'h5 : 3'h0; // @[Fetch.scala 95:39]
  wire [2:0] _T_15 = 4'h2 == _T_5 ? 3'h1 : waiting; // @[Mux.scala 81:58]
  wire [2:0] _T_17 = 4'h4 == _T_5 ? 3'h2 : _T_15; // @[Mux.scala 81:58]
  wire [2:0] _T_19 = 4'h5 == _T_5 ? 3'h3 : _T_17; // @[Mux.scala 81:58]
  wire [2:0] _T_21 = 4'h6 == _T_5 ? 3'h4 : _T_19; // @[Mux.scala 81:58]
  wire [2:0] _T_23 = 4'h3 == _T_5 ? _T_12 : _T_21; // @[Mux.scala 81:58]
  wire [2:0] _T_25 = 4'h7 == _T_5 ? 3'h6 : _T_23; // @[Mux.scala 81:58]
  wire [2:0] nextWait = _T_4 ? waiting : _T_25; // @[Fetch.scala 84:19]
  wire  _T_29 = _T_1 | ~io_fetchBuffer_toBuffer_0_valid; // @[Fetch.scala 108:25]
  wire  _T_30 = checkBranches_0_io_branchType == 4'h3; // @[Fetch.scala 109:31]
  wire  _T_31 = checkBranches_0_io_branchType == 4'h2; // @[Fetch.scala 110:31]
  wire  _T_32 = nextWait != 3'h0; // @[Fetch.scala 111:19]
  wire  _T_33 = checkBranches_0_io_branchType == 4'h1; // @[Fetch.scala 112:31]
  wire [3:0] _T_34 = _T_33 ? $signed(4'sh2) : $signed(4'sh4); // @[Mux.scala 101:16]
  wire [3:0] _T_35 = _T_32 ? $signed(4'sh0) : $signed(_T_34); // @[Mux.scala 101:16]
  wire [3:0] _T_36 = _T_31 ? $signed(4'sh0) : $signed(_T_35); // @[Mux.scala 101:16]
  wire [20:0] _T_37 = _T_30 ? $signed(checkBranches_0_io_offset) : $signed({{17{_T_36[3]}},_T_36}); // @[Mux.scala 101:16]
  wire [20:0] _T_38 = _T_29 ? $signed(21'sh0) : $signed(_T_37); // @[Mux.scala 101:16]
  wire [63:0] _GEN_21 = {{43{_T_38[20]}},_T_38}; // @[Fetch.scala 105:29]
  wire [63:0] nextPC = $signed(pc) + $signed(_GEN_21); // @[Fetch.scala 114:8]
  wire [63:0] _pc_T_4 = $signed(pc) + $signed(io_collectedBranchAddresses_addresses_bits_programCounterOffset); // @[Fetch.scala 125:57]
  wire [2:0] _GEN_0 = io_collectedBranchAddresses_addresses_valid & ~io_collectedBranchAddresses_addresses_bits_threadId
     ? 3'h0 : nextWait; // @[Fetch.scala 117:11 123:55 124:17]
  wire [63:0] _GEN_1 = io_collectedBranchAddresses_addresses_valid & ~
    io_collectedBranchAddresses_addresses_bits_threadId ? _pc_T_4 : nextPC; // @[Fetch.scala 123:55 125:12 116:6]
  wire [2:0] _GEN_2 = waiting == 3'h1 | waiting == 3'h2 ? _GEN_0 : nextWait; // @[Fetch.scala 117:11 121:78]
  wire [63:0] _GEN_3 = waiting == 3'h1 | waiting == 3'h2 ? _GEN_1 : nextPC; // @[Fetch.scala 116:6 121:78]
  wire  _T_52 = io_reorderBufferEmpty & io_loadStoreQueueEmpty & io_fetchBuffer_empty; // @[Fetch.scala 130:57]
  wire [63:0] _pc_T_6 = pc + 64'h4; // @[Fetch.scala 133:18]
  wire [2:0] _GEN_4 = _T_52 ? 3'h0 : _GEN_2; // @[Fetch.scala 131:9 132:17]
  wire [63:0] _GEN_5 = _T_52 ? _pc_T_6 : _GEN_3; // @[Fetch.scala 131:9 133:12]
  wire [2:0] _GEN_6 = waiting == 3'h3 | waiting == 3'h4 ? _GEN_4 : _GEN_2; // @[Fetch.scala 128:79]
  wire [63:0] _GEN_7 = waiting == 3'h3 | waiting == 3'h4 ? _GEN_5 : _GEN_3; // @[Fetch.scala 128:79]
  wire [2:0] _GEN_8 = io_csrReservationStationEmpty ? 3'h0 : _GEN_6; // @[Fetch.scala 142:43 143:17]
  wire [63:0] _GEN_9 = io_csrReservationStationEmpty ? io_csr_mepc : _GEN_7; // @[Fetch.scala 142:43 144:12]
  wire [2:0] _GEN_10 = waiting == 3'h6 ? _GEN_8 : _GEN_6; // @[Fetch.scala 141:42]
  wire [63:0] _GEN_11 = waiting == 3'h6 ? _GEN_9 : _GEN_7; // @[Fetch.scala 141:42]
  wire [63:0] _pc_T_8 = {io_csr_mtvec[63:2],2'h0}; // @[Fetch.scala 151:37]
  wire [62:0] _GEN_22 = {{1'd0}, io_csr_mtvec[63:2]}; // @[Fetch.scala 153:38]
  wire [62:0] _pc_T_12 = _GEN_22 + io_csr_mcause[62:0]; // @[Fetch.scala 153:38]
  wire [64:0] _pc_T_13 = {_pc_T_12,2'h0}; // @[Fetch.scala 153:62]
  wire [64:0] _GEN_12 = io_csr_mcause[1:0] == 2'h1 ? _pc_T_13 : {{1'd0}, _GEN_11}; // @[Fetch.scala 152:49 153:14]
  wire [64:0] _GEN_13 = io_csr_mcause[1:0] == 2'h0 ? {{1'd0}, _pc_T_8} : _GEN_12; // @[Fetch.scala 150:43 151:14]
  wire [2:0] _GEN_14 = io_csrReservationStationEmpty ? 3'h0 : _GEN_10; // @[Fetch.scala 148:43 149:17]
  wire [64:0] _GEN_15 = io_csrReservationStationEmpty ? _GEN_13 : {{1'd0}, _GEN_11}; // @[Fetch.scala 148:43]
  wire [64:0] _GEN_17 = waiting == 3'h7 ? _GEN_15 : {{1'd0}, _GEN_11}; // @[Fetch.scala 147:47]
  wire [64:0] _GEN_19 = _T ? _GEN_17 : {{1'd0}, nextPC}; // @[Fetch.scala 120:40 116:6]
  wire [64:0] _GEN_23 = reset ? 65'h20000000 : _GEN_19; // @[Fetch.scala 57:{19,19}]
  CheckBranch checkBranches_0 ( // @[Fetch.scala 54:63]
    .io_instruction(checkBranches_0_io_instruction),
    .io_branchType(checkBranches_0_io_branchType),
    .io_offset(checkBranches_0_io_offset)
  );
  assign io_cache_0_address_valid = waiting == 3'h0; // @[Fetch.scala 81:37]
  assign io_cache_0_address_bits = pc; // @[Fetch.scala 68:24]
  assign io_fetchBuffer_toBuffer_0_valid = instructionValid & checkBranches_0_io_branchType != 4'h7 & ~io_isError; // @[Fetch.scala 77:83]
  assign io_fetchBuffer_toBuffer_0_bits_instruction = io_cache_0_output_bits; // @[Fetch.scala 79:30]
  assign io_fetchBuffer_toBuffer_0_bits_programCounter = pc; // @[Fetch.scala 78:33]
  assign checkBranches_0_io_instruction = io_cache_0_output_bits; // @[Fetch.scala 71:27]
  always @(posedge clock) begin
    pc <= _GEN_23[63:0]; // @[Fetch.scala 57:{19,19}]
    if (reset) begin // @[Fetch.scala 60:24]
      waiting <= 3'h0; // @[Fetch.scala 60:24]
    end else if (io_isError) begin // @[Fetch.scala 159:20]
      waiting <= 3'h7; // @[Fetch.scala 160:13]
    end else if (_T) begin // @[Fetch.scala 120:40]
      if (waiting == 3'h7) begin // @[Fetch.scala 147:47]
        waiting <= _GEN_14;
      end else begin
        waiting <= _GEN_10;
      end
    end else if (!(_T_4)) begin // @[Fetch.scala 84:19]
      waiting <= _T_25;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  pc = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  waiting = _RAND_1[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Fetch_1(
  input         clock,
  input         reset,
  output        io_cache_0_address_valid,
  output [63:0] io_cache_0_address_bits,
  input         io_cache_0_output_valid,
  input  [31:0] io_cache_0_output_bits,
  input         io_reorderBufferEmpty,
  input         io_loadStoreQueueEmpty,
  input         io_collectedBranchAddresses_addresses_valid,
  input         io_collectedBranchAddresses_addresses_bits_threadId,
  input  [63:0] io_collectedBranchAddresses_addresses_bits_programCounterOffset,
  input         io_fetchBuffer_toBuffer_0_ready,
  output        io_fetchBuffer_toBuffer_0_valid,
  output [31:0] io_fetchBuffer_toBuffer_0_bits_instruction,
  output [63:0] io_fetchBuffer_toBuffer_0_bits_programCounter,
  input         io_fetchBuffer_empty,
  input  [63:0] io_csr_mtvec,
  input  [63:0] io_csr_mepc,
  input  [63:0] io_csr_mcause,
  input         io_csrReservationStationEmpty,
  input         io_isError
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] checkBranches_0_io_instruction; // @[Fetch.scala 54:63]
  wire [3:0] checkBranches_0_io_branchType; // @[Fetch.scala 54:63]
  wire [20:0] checkBranches_0_io_offset; // @[Fetch.scala 54:63]
  reg [63:0] pc; // @[Fetch.scala 57:19]
  reg [2:0] waiting; // @[Fetch.scala 60:24]
  wire  instructionValid = io_cache_0_output_valid & waiting == 3'h0; // @[Fetch.scala 76:47]
  wire  _T = waiting != 3'h0; // @[Fetch.scala 85:16]
  wire  _T_1 = ~io_fetchBuffer_toBuffer_0_ready; // @[Fetch.scala 85:42]
  wire  _T_4 = waiting != 3'h0 | ~io_fetchBuffer_toBuffer_0_ready | ~instructionValid; // @[Fetch.scala 85:57]
  wire [3:0] _T_5 = checkBranches_0_io_branchType; // @[Fetch.scala 88:30]
  wire  _T_11 = $signed(checkBranches_0_io_offset) == 21'sh0; // @[Fetch.scala 96:30]
  wire [2:0] _T_12 = _T_11 ? 3'h5 : 3'h0; // @[Fetch.scala 95:39]
  wire [2:0] _T_15 = 4'h2 == _T_5 ? 3'h1 : waiting; // @[Mux.scala 81:58]
  wire [2:0] _T_17 = 4'h4 == _T_5 ? 3'h2 : _T_15; // @[Mux.scala 81:58]
  wire [2:0] _T_19 = 4'h5 == _T_5 ? 3'h3 : _T_17; // @[Mux.scala 81:58]
  wire [2:0] _T_21 = 4'h6 == _T_5 ? 3'h4 : _T_19; // @[Mux.scala 81:58]
  wire [2:0] _T_23 = 4'h3 == _T_5 ? _T_12 : _T_21; // @[Mux.scala 81:58]
  wire [2:0] _T_25 = 4'h7 == _T_5 ? 3'h6 : _T_23; // @[Mux.scala 81:58]
  wire [2:0] nextWait = _T_4 ? waiting : _T_25; // @[Fetch.scala 84:19]
  wire  _T_29 = _T_1 | ~io_fetchBuffer_toBuffer_0_valid; // @[Fetch.scala 108:25]
  wire  _T_30 = checkBranches_0_io_branchType == 4'h3; // @[Fetch.scala 109:31]
  wire  _T_31 = checkBranches_0_io_branchType == 4'h2; // @[Fetch.scala 110:31]
  wire  _T_32 = nextWait != 3'h0; // @[Fetch.scala 111:19]
  wire  _T_33 = checkBranches_0_io_branchType == 4'h1; // @[Fetch.scala 112:31]
  wire [3:0] _T_34 = _T_33 ? $signed(4'sh2) : $signed(4'sh4); // @[Mux.scala 101:16]
  wire [3:0] _T_35 = _T_32 ? $signed(4'sh0) : $signed(_T_34); // @[Mux.scala 101:16]
  wire [3:0] _T_36 = _T_31 ? $signed(4'sh0) : $signed(_T_35); // @[Mux.scala 101:16]
  wire [20:0] _T_37 = _T_30 ? $signed(checkBranches_0_io_offset) : $signed({{17{_T_36[3]}},_T_36}); // @[Mux.scala 101:16]
  wire [20:0] _T_38 = _T_29 ? $signed(21'sh0) : $signed(_T_37); // @[Mux.scala 101:16]
  wire [63:0] _GEN_21 = {{43{_T_38[20]}},_T_38}; // @[Fetch.scala 105:29]
  wire [63:0] nextPC = $signed(pc) + $signed(_GEN_21); // @[Fetch.scala 114:8]
  wire [63:0] _pc_T_4 = $signed(pc) + $signed(io_collectedBranchAddresses_addresses_bits_programCounterOffset); // @[Fetch.scala 125:57]
  wire [2:0] _GEN_0 = io_collectedBranchAddresses_addresses_valid & io_collectedBranchAddresses_addresses_bits_threadId
     ? 3'h0 : nextWait; // @[Fetch.scala 117:11 123:55 124:17]
  wire [63:0] _GEN_1 = io_collectedBranchAddresses_addresses_valid & io_collectedBranchAddresses_addresses_bits_threadId
     ? _pc_T_4 : nextPC; // @[Fetch.scala 123:55 125:12 116:6]
  wire [2:0] _GEN_2 = waiting == 3'h1 | waiting == 3'h2 ? _GEN_0 : nextWait; // @[Fetch.scala 117:11 121:78]
  wire [63:0] _GEN_3 = waiting == 3'h1 | waiting == 3'h2 ? _GEN_1 : nextPC; // @[Fetch.scala 116:6 121:78]
  wire  _T_52 = io_reorderBufferEmpty & io_loadStoreQueueEmpty & io_fetchBuffer_empty; // @[Fetch.scala 130:57]
  wire [63:0] _pc_T_6 = pc + 64'h4; // @[Fetch.scala 133:18]
  wire [2:0] _GEN_4 = _T_52 ? 3'h0 : _GEN_2; // @[Fetch.scala 131:9 132:17]
  wire [63:0] _GEN_5 = _T_52 ? _pc_T_6 : _GEN_3; // @[Fetch.scala 131:9 133:12]
  wire [2:0] _GEN_6 = waiting == 3'h3 | waiting == 3'h4 ? _GEN_4 : _GEN_2; // @[Fetch.scala 128:79]
  wire [63:0] _GEN_7 = waiting == 3'h3 | waiting == 3'h4 ? _GEN_5 : _GEN_3; // @[Fetch.scala 128:79]
  wire [2:0] _GEN_8 = io_csrReservationStationEmpty ? 3'h0 : _GEN_6; // @[Fetch.scala 142:43 143:17]
  wire [63:0] _GEN_9 = io_csrReservationStationEmpty ? io_csr_mepc : _GEN_7; // @[Fetch.scala 142:43 144:12]
  wire [2:0] _GEN_10 = waiting == 3'h6 ? _GEN_8 : _GEN_6; // @[Fetch.scala 141:42]
  wire [63:0] _GEN_11 = waiting == 3'h6 ? _GEN_9 : _GEN_7; // @[Fetch.scala 141:42]
  wire [63:0] _pc_T_8 = {io_csr_mtvec[63:2],2'h0}; // @[Fetch.scala 151:37]
  wire [62:0] _GEN_22 = {{1'd0}, io_csr_mtvec[63:2]}; // @[Fetch.scala 153:38]
  wire [62:0] _pc_T_12 = _GEN_22 + io_csr_mcause[62:0]; // @[Fetch.scala 153:38]
  wire [64:0] _pc_T_13 = {_pc_T_12,2'h0}; // @[Fetch.scala 153:62]
  wire [64:0] _GEN_12 = io_csr_mcause[1:0] == 2'h1 ? _pc_T_13 : {{1'd0}, _GEN_11}; // @[Fetch.scala 152:49 153:14]
  wire [64:0] _GEN_13 = io_csr_mcause[1:0] == 2'h0 ? {{1'd0}, _pc_T_8} : _GEN_12; // @[Fetch.scala 150:43 151:14]
  wire [2:0] _GEN_14 = io_csrReservationStationEmpty ? 3'h0 : _GEN_10; // @[Fetch.scala 148:43 149:17]
  wire [64:0] _GEN_15 = io_csrReservationStationEmpty ? _GEN_13 : {{1'd0}, _GEN_11}; // @[Fetch.scala 148:43]
  wire [64:0] _GEN_17 = waiting == 3'h7 ? _GEN_15 : {{1'd0}, _GEN_11}; // @[Fetch.scala 147:47]
  wire [64:0] _GEN_19 = _T ? _GEN_17 : {{1'd0}, nextPC}; // @[Fetch.scala 120:40 116:6]
  wire [64:0] _GEN_23 = reset ? 65'h20000000 : _GEN_19; // @[Fetch.scala 57:{19,19}]
  CheckBranch checkBranches_0 ( // @[Fetch.scala 54:63]
    .io_instruction(checkBranches_0_io_instruction),
    .io_branchType(checkBranches_0_io_branchType),
    .io_offset(checkBranches_0_io_offset)
  );
  assign io_cache_0_address_valid = waiting == 3'h0; // @[Fetch.scala 81:37]
  assign io_cache_0_address_bits = pc; // @[Fetch.scala 68:24]
  assign io_fetchBuffer_toBuffer_0_valid = instructionValid & checkBranches_0_io_branchType != 4'h7 & ~io_isError; // @[Fetch.scala 77:83]
  assign io_fetchBuffer_toBuffer_0_bits_instruction = io_cache_0_output_bits; // @[Fetch.scala 79:30]
  assign io_fetchBuffer_toBuffer_0_bits_programCounter = pc; // @[Fetch.scala 78:33]
  assign checkBranches_0_io_instruction = io_cache_0_output_bits; // @[Fetch.scala 71:27]
  always @(posedge clock) begin
    pc <= _GEN_23[63:0]; // @[Fetch.scala 57:{19,19}]
    if (reset) begin // @[Fetch.scala 60:24]
      waiting <= 3'h0; // @[Fetch.scala 60:24]
    end else if (io_isError) begin // @[Fetch.scala 159:20]
      waiting <= 3'h7; // @[Fetch.scala 160:13]
    end else if (_T) begin // @[Fetch.scala 120:40]
      if (waiting == 3'h7) begin // @[Fetch.scala 147:47]
        waiting <= _GEN_14;
      end else begin
        waiting <= _GEN_10;
      end
    end else if (!(_T_4)) begin // @[Fetch.scala 84:19]
      waiting <= _T_25;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  pc = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  waiting = _RAND_1[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module FetchBuffer(
  input         clock,
  input         reset,
  input         io_output_0_ready,
  output        io_output_0_valid,
  output [31:0] io_output_0_bits_instruction,
  output [63:0] io_output_0_bits_programCounter,
  output        io_input_toBuffer_0_ready,
  input         io_input_toBuffer_0_valid,
  input  [31:0] io_input_toBuffer_0_bits_instruction,
  input  [63:0] io_input_toBuffer_0_bits_programCounter,
  output        io_input_empty
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] buffer_0_instruction; // @[FetchBuffer.scala 16:19]
  reg [63:0] buffer_0_programCounter; // @[FetchBuffer.scala 16:19]
  reg [31:0] buffer_1_instruction; // @[FetchBuffer.scala 16:19]
  reg [63:0] buffer_1_programCounter; // @[FetchBuffer.scala 16:19]
  reg [31:0] buffer_2_instruction; // @[FetchBuffer.scala 16:19]
  reg [63:0] buffer_2_programCounter; // @[FetchBuffer.scala 16:19]
  reg [31:0] buffer_3_instruction; // @[FetchBuffer.scala 16:19]
  reg [63:0] buffer_3_programCounter; // @[FetchBuffer.scala 16:19]
  reg [1:0] head; // @[FetchBuffer.scala 20:21]
  reg [1:0] tail; // @[FetchBuffer.scala 21:21]
  wire [1:0] _indexOk_T_1 = head + 2'h1; // @[FetchBuffer.scala 27:30]
  wire  indexOk = _indexOk_T_1 != tail; // @[FetchBuffer.scala 27:36]
  wire  valid = io_input_toBuffer_0_valid & indexOk; // @[FetchBuffer.scala 29:27]
  wire  indexOk_1 = tail != head; // @[FetchBuffer.scala 44:30]
  wire  valid_1 = io_output_0_ready & indexOk_1; // @[FetchBuffer.scala 46:27]
  wire [31:0] _GEN_17 = 2'h1 == tail ? buffer_1_instruction : buffer_0_instruction; // @[FetchBuffer.scala 50:{28,28}]
  wire [31:0] _GEN_18 = 2'h2 == tail ? buffer_2_instruction : _GEN_17; // @[FetchBuffer.scala 50:{28,28}]
  wire [31:0] _GEN_19 = 2'h3 == tail ? buffer_3_instruction : _GEN_18; // @[FetchBuffer.scala 50:{28,28}]
  wire [63:0] _GEN_21 = 2'h1 == tail ? buffer_1_programCounter : buffer_0_programCounter; // @[FetchBuffer.scala 51:{31,31}]
  wire [63:0] _GEN_22 = 2'h2 == tail ? buffer_2_programCounter : _GEN_21; // @[FetchBuffer.scala 51:{31,31}]
  wire [63:0] _GEN_23 = 2'h3 == tail ? buffer_3_programCounter : _GEN_22; // @[FetchBuffer.scala 51:{31,31}]
  wire [1:0] _T_4 = tail + 2'h1; // @[FetchBuffer.scala 53:38]
  assign io_output_0_valid = tail != head; // @[FetchBuffer.scala 44:30]
  assign io_output_0_bits_instruction = valid_1 ? _GEN_19 : 32'h0; // @[FetchBuffer.scala 49:19 47:26 50:28]
  assign io_output_0_bits_programCounter = valid_1 ? _GEN_23 : 64'h0; // @[FetchBuffer.scala 49:19 48:29 51:31]
  assign io_input_toBuffer_0_ready = _indexOk_T_1 != tail; // @[FetchBuffer.scala 27:36]
  assign io_input_empty = head == tail; // @[FetchBuffer.scala 22:26]
  always @(posedge clock) begin
    if (valid) begin // @[FetchBuffer.scala 30:19]
      if (2'h0 == head) begin // @[FetchBuffer.scala 31:26]
        buffer_0_instruction <= io_input_toBuffer_0_bits_instruction; // @[FetchBuffer.scala 31:26]
      end
    end
    if (valid) begin // @[FetchBuffer.scala 30:19]
      if (2'h0 == head) begin // @[FetchBuffer.scala 31:26]
        buffer_0_programCounter <= io_input_toBuffer_0_bits_programCounter; // @[FetchBuffer.scala 31:26]
      end
    end
    if (valid) begin // @[FetchBuffer.scala 30:19]
      if (2'h1 == head) begin // @[FetchBuffer.scala 31:26]
        buffer_1_instruction <= io_input_toBuffer_0_bits_instruction; // @[FetchBuffer.scala 31:26]
      end
    end
    if (valid) begin // @[FetchBuffer.scala 30:19]
      if (2'h1 == head) begin // @[FetchBuffer.scala 31:26]
        buffer_1_programCounter <= io_input_toBuffer_0_bits_programCounter; // @[FetchBuffer.scala 31:26]
      end
    end
    if (valid) begin // @[FetchBuffer.scala 30:19]
      if (2'h2 == head) begin // @[FetchBuffer.scala 31:26]
        buffer_2_instruction <= io_input_toBuffer_0_bits_instruction; // @[FetchBuffer.scala 31:26]
      end
    end
    if (valid) begin // @[FetchBuffer.scala 30:19]
      if (2'h2 == head) begin // @[FetchBuffer.scala 31:26]
        buffer_2_programCounter <= io_input_toBuffer_0_bits_programCounter; // @[FetchBuffer.scala 31:26]
      end
    end
    if (valid) begin // @[FetchBuffer.scala 30:19]
      if (2'h3 == head) begin // @[FetchBuffer.scala 31:26]
        buffer_3_instruction <= io_input_toBuffer_0_bits_instruction; // @[FetchBuffer.scala 31:26]
      end
    end
    if (valid) begin // @[FetchBuffer.scala 30:19]
      if (2'h3 == head) begin // @[FetchBuffer.scala 31:26]
        buffer_3_programCounter <= io_input_toBuffer_0_bits_programCounter; // @[FetchBuffer.scala 31:26]
      end
    end
    if (reset) begin // @[FetchBuffer.scala 20:21]
      head <= 2'h0; // @[FetchBuffer.scala 20:21]
    end else if (valid) begin // @[FetchBuffer.scala 36:21]
      head <= _indexOk_T_1;
    end
    if (reset) begin // @[FetchBuffer.scala 21:21]
      tail <= 2'h0; // @[FetchBuffer.scala 21:21]
    end else if (valid_1) begin // @[FetchBuffer.scala 53:21]
      tail <= _T_4;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  buffer_0_instruction = _RAND_0[31:0];
  _RAND_1 = {2{`RANDOM}};
  buffer_0_programCounter = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  buffer_1_instruction = _RAND_2[31:0];
  _RAND_3 = {2{`RANDOM}};
  buffer_1_programCounter = _RAND_3[63:0];
  _RAND_4 = {1{`RANDOM}};
  buffer_2_instruction = _RAND_4[31:0];
  _RAND_5 = {2{`RANDOM}};
  buffer_2_programCounter = _RAND_5[63:0];
  _RAND_6 = {1{`RANDOM}};
  buffer_3_instruction = _RAND_6[31:0];
  _RAND_7 = {2{`RANDOM}};
  buffer_3_programCounter = _RAND_7[63:0];
  _RAND_8 = {1{`RANDOM}};
  head = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  tail = _RAND_9[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ReorderBuffer(
  input         clock,
  input         reset,
  input  [4:0]  io_decoders_0_source1_sourceRegister,
  output        io_decoders_0_source1_matchingTag_valid,
  output [3:0]  io_decoders_0_source1_matchingTag_bits_id,
  output        io_decoders_0_source1_value_valid,
  output [63:0] io_decoders_0_source1_value_bits,
  input  [4:0]  io_decoders_0_source2_sourceRegister,
  output        io_decoders_0_source2_matchingTag_valid,
  output [3:0]  io_decoders_0_source2_matchingTag_bits_id,
  output        io_decoders_0_source2_value_valid,
  output [63:0] io_decoders_0_source2_value_bits,
  input  [4:0]  io_decoders_0_destination_destinationRegister,
  output [3:0]  io_decoders_0_destination_destinationTag_id,
  input         io_decoders_0_destination_storeSign,
  output        io_decoders_0_ready,
  input         io_decoders_0_valid,
  input         io_collectedOutputs_outputs_valid,
  input         io_collectedOutputs_outputs_bits_resultType,
  input  [63:0] io_collectedOutputs_outputs_bits_value,
  input         io_collectedOutputs_outputs_bits_isError,
  input         io_collectedOutputs_outputs_bits_tag_threadId,
  input  [3:0]  io_collectedOutputs_outputs_bits_tag_id,
  output        io_registerFile_0_valid,
  output [4:0]  io_registerFile_0_bits_destinationRegister,
  output [63:0] io_registerFile_0_bits_value,
  output        io_registerFile_1_valid,
  output [4:0]  io_registerFile_1_bits_destinationRegister,
  output [63:0] io_registerFile_1_bits_value,
  output        io_registerFile_2_valid,
  output [4:0]  io_registerFile_2_bits_destinationRegister,
  output [63:0] io_registerFile_2_bits_value,
  output        io_registerFile_3_valid,
  output [4:0]  io_registerFile_3_bits_destinationRegister,
  output [63:0] io_registerFile_3_bits_value,
  output        io_loadStoreQueue_0_valid,
  output [3:0]  io_loadStoreQueue_0_bits_destinationTag_id,
  output        io_loadStoreQueue_1_valid,
  output [3:0]  io_loadStoreQueue_1_bits_destinationTag_id,
  output        io_loadStoreQueue_2_valid,
  output [3:0]  io_loadStoreQueue_2_bits_destinationTag_id,
  output        io_loadStoreQueue_3_valid,
  output [3:0]  io_loadStoreQueue_3_bits_destinationTag_id,
  output        io_isEmpty,
  output [1:0]  io_csr_retireCount,
  output        io_isError
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [63:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [63:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [63:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [63:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [63:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [63:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [63:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [63:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] head; // @[ReorderBuffer.scala 53:21]
  reg [3:0] tail; // @[ReorderBuffer.scala 54:21]
  reg [4:0] buffer_0_destinationRegister; // @[ReorderBuffer.scala 55:23]
  reg  buffer_0_valueReady; // @[ReorderBuffer.scala 55:23]
  reg [63:0] buffer_0_value; // @[ReorderBuffer.scala 55:23]
  reg  buffer_0_storeSign; // @[ReorderBuffer.scala 55:23]
  reg  buffer_0_isError; // @[ReorderBuffer.scala 55:23]
  reg [4:0] buffer_1_destinationRegister; // @[ReorderBuffer.scala 55:23]
  reg  buffer_1_valueReady; // @[ReorderBuffer.scala 55:23]
  reg [63:0] buffer_1_value; // @[ReorderBuffer.scala 55:23]
  reg  buffer_1_storeSign; // @[ReorderBuffer.scala 55:23]
  reg  buffer_1_isError; // @[ReorderBuffer.scala 55:23]
  reg [4:0] buffer_2_destinationRegister; // @[ReorderBuffer.scala 55:23]
  reg  buffer_2_valueReady; // @[ReorderBuffer.scala 55:23]
  reg [63:0] buffer_2_value; // @[ReorderBuffer.scala 55:23]
  reg  buffer_2_storeSign; // @[ReorderBuffer.scala 55:23]
  reg  buffer_2_isError; // @[ReorderBuffer.scala 55:23]
  reg [4:0] buffer_3_destinationRegister; // @[ReorderBuffer.scala 55:23]
  reg  buffer_3_valueReady; // @[ReorderBuffer.scala 55:23]
  reg [63:0] buffer_3_value; // @[ReorderBuffer.scala 55:23]
  reg  buffer_3_storeSign; // @[ReorderBuffer.scala 55:23]
  reg  buffer_3_isError; // @[ReorderBuffer.scala 55:23]
  reg [4:0] buffer_4_destinationRegister; // @[ReorderBuffer.scala 55:23]
  reg  buffer_4_valueReady; // @[ReorderBuffer.scala 55:23]
  reg [63:0] buffer_4_value; // @[ReorderBuffer.scala 55:23]
  reg  buffer_4_storeSign; // @[ReorderBuffer.scala 55:23]
  reg  buffer_4_isError; // @[ReorderBuffer.scala 55:23]
  reg [4:0] buffer_5_destinationRegister; // @[ReorderBuffer.scala 55:23]
  reg  buffer_5_valueReady; // @[ReorderBuffer.scala 55:23]
  reg [63:0] buffer_5_value; // @[ReorderBuffer.scala 55:23]
  reg  buffer_5_storeSign; // @[ReorderBuffer.scala 55:23]
  reg  buffer_5_isError; // @[ReorderBuffer.scala 55:23]
  reg [4:0] buffer_6_destinationRegister; // @[ReorderBuffer.scala 55:23]
  reg  buffer_6_valueReady; // @[ReorderBuffer.scala 55:23]
  reg [63:0] buffer_6_value; // @[ReorderBuffer.scala 55:23]
  reg  buffer_6_storeSign; // @[ReorderBuffer.scala 55:23]
  reg  buffer_6_isError; // @[ReorderBuffer.scala 55:23]
  reg [4:0] buffer_7_destinationRegister; // @[ReorderBuffer.scala 55:23]
  reg  buffer_7_valueReady; // @[ReorderBuffer.scala 55:23]
  reg [63:0] buffer_7_value; // @[ReorderBuffer.scala 55:23]
  reg  buffer_7_storeSign; // @[ReorderBuffer.scala 55:23]
  reg  buffer_7_isError; // @[ReorderBuffer.scala 55:23]
  reg [4:0] buffer_8_destinationRegister; // @[ReorderBuffer.scala 55:23]
  reg  buffer_8_valueReady; // @[ReorderBuffer.scala 55:23]
  reg [63:0] buffer_8_value; // @[ReorderBuffer.scala 55:23]
  reg  buffer_8_storeSign; // @[ReorderBuffer.scala 55:23]
  reg  buffer_8_isError; // @[ReorderBuffer.scala 55:23]
  reg [4:0] buffer_9_destinationRegister; // @[ReorderBuffer.scala 55:23]
  reg  buffer_9_valueReady; // @[ReorderBuffer.scala 55:23]
  reg [63:0] buffer_9_value; // @[ReorderBuffer.scala 55:23]
  reg  buffer_9_storeSign; // @[ReorderBuffer.scala 55:23]
  reg  buffer_9_isError; // @[ReorderBuffer.scala 55:23]
  reg [4:0] buffer_10_destinationRegister; // @[ReorderBuffer.scala 55:23]
  reg  buffer_10_valueReady; // @[ReorderBuffer.scala 55:23]
  reg [63:0] buffer_10_value; // @[ReorderBuffer.scala 55:23]
  reg  buffer_10_storeSign; // @[ReorderBuffer.scala 55:23]
  reg  buffer_10_isError; // @[ReorderBuffer.scala 55:23]
  reg [4:0] buffer_11_destinationRegister; // @[ReorderBuffer.scala 55:23]
  reg  buffer_11_valueReady; // @[ReorderBuffer.scala 55:23]
  reg [63:0] buffer_11_value; // @[ReorderBuffer.scala 55:23]
  reg  buffer_11_storeSign; // @[ReorderBuffer.scala 55:23]
  reg  buffer_11_isError; // @[ReorderBuffer.scala 55:23]
  reg [4:0] buffer_12_destinationRegister; // @[ReorderBuffer.scala 55:23]
  reg  buffer_12_valueReady; // @[ReorderBuffer.scala 55:23]
  reg [63:0] buffer_12_value; // @[ReorderBuffer.scala 55:23]
  reg  buffer_12_storeSign; // @[ReorderBuffer.scala 55:23]
  reg  buffer_12_isError; // @[ReorderBuffer.scala 55:23]
  reg [4:0] buffer_13_destinationRegister; // @[ReorderBuffer.scala 55:23]
  reg  buffer_13_valueReady; // @[ReorderBuffer.scala 55:23]
  reg [63:0] buffer_13_value; // @[ReorderBuffer.scala 55:23]
  reg  buffer_13_storeSign; // @[ReorderBuffer.scala 55:23]
  reg  buffer_13_isError; // @[ReorderBuffer.scala 55:23]
  reg [4:0] buffer_14_destinationRegister; // @[ReorderBuffer.scala 55:23]
  reg  buffer_14_valueReady; // @[ReorderBuffer.scala 55:23]
  reg [63:0] buffer_14_value; // @[ReorderBuffer.scala 55:23]
  reg  buffer_14_storeSign; // @[ReorderBuffer.scala 55:23]
  reg  buffer_14_isError; // @[ReorderBuffer.scala 55:23]
  reg [4:0] buffer_15_destinationRegister; // @[ReorderBuffer.scala 55:23]
  reg  buffer_15_valueReady; // @[ReorderBuffer.scala 55:23]
  reg [63:0] buffer_15_value; // @[ReorderBuffer.scala 55:23]
  reg  buffer_15_storeSign; // @[ReorderBuffer.scala 55:23]
  reg  buffer_15_isError; // @[ReorderBuffer.scala 55:23]
  reg  registerTagMap_1_valid; // @[ReorderBuffer.scala 69:39]
  reg [3:0] registerTagMap_1_tagId; // @[ReorderBuffer.scala 69:39]
  reg  registerTagMap_2_valid; // @[ReorderBuffer.scala 69:39]
  reg [3:0] registerTagMap_2_tagId; // @[ReorderBuffer.scala 69:39]
  reg  registerTagMap_3_valid; // @[ReorderBuffer.scala 69:39]
  reg [3:0] registerTagMap_3_tagId; // @[ReorderBuffer.scala 69:39]
  reg  registerTagMap_4_valid; // @[ReorderBuffer.scala 69:39]
  reg [3:0] registerTagMap_4_tagId; // @[ReorderBuffer.scala 69:39]
  reg  registerTagMap_5_valid; // @[ReorderBuffer.scala 69:39]
  reg [3:0] registerTagMap_5_tagId; // @[ReorderBuffer.scala 69:39]
  reg  registerTagMap_6_valid; // @[ReorderBuffer.scala 69:39]
  reg [3:0] registerTagMap_6_tagId; // @[ReorderBuffer.scala 69:39]
  reg  registerTagMap_7_valid; // @[ReorderBuffer.scala 69:39]
  reg [3:0] registerTagMap_7_tagId; // @[ReorderBuffer.scala 69:39]
  reg  registerTagMap_8_valid; // @[ReorderBuffer.scala 69:39]
  reg [3:0] registerTagMap_8_tagId; // @[ReorderBuffer.scala 69:39]
  reg  registerTagMap_9_valid; // @[ReorderBuffer.scala 69:39]
  reg [3:0] registerTagMap_9_tagId; // @[ReorderBuffer.scala 69:39]
  reg  registerTagMap_10_valid; // @[ReorderBuffer.scala 69:39]
  reg [3:0] registerTagMap_10_tagId; // @[ReorderBuffer.scala 69:39]
  reg  registerTagMap_11_valid; // @[ReorderBuffer.scala 69:39]
  reg [3:0] registerTagMap_11_tagId; // @[ReorderBuffer.scala 69:39]
  reg  registerTagMap_12_valid; // @[ReorderBuffer.scala 69:39]
  reg [3:0] registerTagMap_12_tagId; // @[ReorderBuffer.scala 69:39]
  reg  registerTagMap_13_valid; // @[ReorderBuffer.scala 69:39]
  reg [3:0] registerTagMap_13_tagId; // @[ReorderBuffer.scala 69:39]
  reg  registerTagMap_14_valid; // @[ReorderBuffer.scala 69:39]
  reg [3:0] registerTagMap_14_tagId; // @[ReorderBuffer.scala 69:39]
  reg  registerTagMap_15_valid; // @[ReorderBuffer.scala 69:39]
  reg [3:0] registerTagMap_15_tagId; // @[ReorderBuffer.scala 69:39]
  reg  registerTagMap_16_valid; // @[ReorderBuffer.scala 69:39]
  reg [3:0] registerTagMap_16_tagId; // @[ReorderBuffer.scala 69:39]
  reg  registerTagMap_17_valid; // @[ReorderBuffer.scala 69:39]
  reg [3:0] registerTagMap_17_tagId; // @[ReorderBuffer.scala 69:39]
  reg  registerTagMap_18_valid; // @[ReorderBuffer.scala 69:39]
  reg [3:0] registerTagMap_18_tagId; // @[ReorderBuffer.scala 69:39]
  reg  registerTagMap_19_valid; // @[ReorderBuffer.scala 69:39]
  reg [3:0] registerTagMap_19_tagId; // @[ReorderBuffer.scala 69:39]
  reg  registerTagMap_20_valid; // @[ReorderBuffer.scala 69:39]
  reg [3:0] registerTagMap_20_tagId; // @[ReorderBuffer.scala 69:39]
  reg  registerTagMap_21_valid; // @[ReorderBuffer.scala 69:39]
  reg [3:0] registerTagMap_21_tagId; // @[ReorderBuffer.scala 69:39]
  reg  registerTagMap_22_valid; // @[ReorderBuffer.scala 69:39]
  reg [3:0] registerTagMap_22_tagId; // @[ReorderBuffer.scala 69:39]
  reg  registerTagMap_23_valid; // @[ReorderBuffer.scala 69:39]
  reg [3:0] registerTagMap_23_tagId; // @[ReorderBuffer.scala 69:39]
  reg  registerTagMap_24_valid; // @[ReorderBuffer.scala 69:39]
  reg [3:0] registerTagMap_24_tagId; // @[ReorderBuffer.scala 69:39]
  reg  registerTagMap_25_valid; // @[ReorderBuffer.scala 69:39]
  reg [3:0] registerTagMap_25_tagId; // @[ReorderBuffer.scala 69:39]
  reg  registerTagMap_26_valid; // @[ReorderBuffer.scala 69:39]
  reg [3:0] registerTagMap_26_tagId; // @[ReorderBuffer.scala 69:39]
  reg  registerTagMap_27_valid; // @[ReorderBuffer.scala 69:39]
  reg [3:0] registerTagMap_27_tagId; // @[ReorderBuffer.scala 69:39]
  reg  registerTagMap_28_valid; // @[ReorderBuffer.scala 69:39]
  reg [3:0] registerTagMap_28_tagId; // @[ReorderBuffer.scala 69:39]
  reg  registerTagMap_29_valid; // @[ReorderBuffer.scala 69:39]
  reg [3:0] registerTagMap_29_tagId; // @[ReorderBuffer.scala 69:39]
  reg  registerTagMap_30_valid; // @[ReorderBuffer.scala 69:39]
  reg [3:0] registerTagMap_30_tagId; // @[ReorderBuffer.scala 69:39]
  reg  registerTagMap_31_valid; // @[ReorderBuffer.scala 69:39]
  reg [3:0] registerTagMap_31_tagId; // @[ReorderBuffer.scala 69:39]
  wire [4:0] _index_T = {{1'd0}, tail}; // @[ReorderBuffer.scala 77:22]
  wire [3:0] index = _index_T[3:0]; // @[ReorderBuffer.scala 77:22]
  wire  _GEN_1 = 4'h1 == index ? buffer_1_valueReady : buffer_0_valueReady; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_2 = 4'h2 == index ? buffer_2_valueReady : _GEN_1; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_3 = 4'h3 == index ? buffer_3_valueReady : _GEN_2; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_4 = 4'h4 == index ? buffer_4_valueReady : _GEN_3; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_5 = 4'h5 == index ? buffer_5_valueReady : _GEN_4; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_6 = 4'h6 == index ? buffer_6_valueReady : _GEN_5; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_7 = 4'h7 == index ? buffer_7_valueReady : _GEN_6; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_8 = 4'h8 == index ? buffer_8_valueReady : _GEN_7; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_9 = 4'h9 == index ? buffer_9_valueReady : _GEN_8; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_10 = 4'ha == index ? buffer_10_valueReady : _GEN_9; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_11 = 4'hb == index ? buffer_11_valueReady : _GEN_10; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_12 = 4'hc == index ? buffer_12_valueReady : _GEN_11; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_13 = 4'hd == index ? buffer_13_valueReady : _GEN_12; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_14 = 4'he == index ? buffer_14_valueReady : _GEN_13; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_15 = 4'hf == index ? buffer_15_valueReady : _GEN_14; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_17 = 4'h1 == index ? buffer_1_storeSign : buffer_0_storeSign; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_18 = 4'h2 == index ? buffer_2_storeSign : _GEN_17; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_19 = 4'h3 == index ? buffer_3_storeSign : _GEN_18; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_20 = 4'h4 == index ? buffer_4_storeSign : _GEN_19; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_21 = 4'h5 == index ? buffer_5_storeSign : _GEN_20; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_22 = 4'h6 == index ? buffer_6_storeSign : _GEN_21; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_23 = 4'h7 == index ? buffer_7_storeSign : _GEN_22; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_24 = 4'h8 == index ? buffer_8_storeSign : _GEN_23; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_25 = 4'h9 == index ? buffer_9_storeSign : _GEN_24; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_26 = 4'ha == index ? buffer_10_storeSign : _GEN_25; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_27 = 4'hb == index ? buffer_11_storeSign : _GEN_26; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_28 = 4'hc == index ? buffer_12_storeSign : _GEN_27; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_29 = 4'hd == index ? buffer_13_storeSign : _GEN_28; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_30 = 4'he == index ? buffer_14_storeSign : _GEN_29; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_31 = 4'hf == index ? buffer_15_storeSign : _GEN_30; // @[ReorderBuffer.scala 79:{50,50}]
  wire  instructionOk = _GEN_15 | _GEN_31; // @[ReorderBuffer.scala 79:50]
  wire  canCommit = index != head & instructionOk; // @[ReorderBuffer.scala 80:49]
  wire  _GEN_33 = 4'h1 == index ? buffer_1_isError : buffer_0_isError; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_34 = 4'h2 == index ? buffer_2_isError : _GEN_33; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_35 = 4'h3 == index ? buffer_3_isError : _GEN_34; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_36 = 4'h4 == index ? buffer_4_isError : _GEN_35; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_37 = 4'h5 == index ? buffer_5_isError : _GEN_36; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_38 = 4'h6 == index ? buffer_6_isError : _GEN_37; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_39 = 4'h7 == index ? buffer_7_isError : _GEN_38; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_40 = 4'h8 == index ? buffer_8_isError : _GEN_39; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_41 = 4'h9 == index ? buffer_9_isError : _GEN_40; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_42 = 4'ha == index ? buffer_10_isError : _GEN_41; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_43 = 4'hb == index ? buffer_11_isError : _GEN_42; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_44 = 4'hc == index ? buffer_12_isError : _GEN_43; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_45 = 4'hd == index ? buffer_13_isError : _GEN_44; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_46 = 4'he == index ? buffer_14_isError : _GEN_45; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_47 = 4'hf == index ? buffer_15_isError : _GEN_46; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _io_registerFile_0_valid_T = ~_GEN_47; // @[ReorderBuffer.scala 83:30]
  wire [63:0] _GEN_49 = 4'h1 == index ? buffer_1_value : buffer_0_value; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_50 = 4'h2 == index ? buffer_2_value : _GEN_49; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_51 = 4'h3 == index ? buffer_3_value : _GEN_50; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_52 = 4'h4 == index ? buffer_4_value : _GEN_51; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_53 = 4'h5 == index ? buffer_5_value : _GEN_52; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_54 = 4'h6 == index ? buffer_6_value : _GEN_53; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_55 = 4'h7 == index ? buffer_7_value : _GEN_54; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_56 = 4'h8 == index ? buffer_8_value : _GEN_55; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_57 = 4'h9 == index ? buffer_9_value : _GEN_56; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_58 = 4'ha == index ? buffer_10_value : _GEN_57; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_59 = 4'hb == index ? buffer_11_value : _GEN_58; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_60 = 4'hc == index ? buffer_12_value : _GEN_59; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_61 = 4'hd == index ? buffer_13_value : _GEN_60; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_62 = 4'he == index ? buffer_14_value : _GEN_61; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_63 = 4'hf == index ? buffer_15_value : _GEN_62; // @[ReorderBuffer.scala 90:{23,23}]
  wire [4:0] _GEN_65 = 4'h1 == index ? buffer_1_destinationRegister : buffer_0_destinationRegister; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_66 = 4'h2 == index ? buffer_2_destinationRegister : _GEN_65; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_67 = 4'h3 == index ? buffer_3_destinationRegister : _GEN_66; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_68 = 4'h4 == index ? buffer_4_destinationRegister : _GEN_67; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_69 = 4'h5 == index ? buffer_5_destinationRegister : _GEN_68; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_70 = 4'h6 == index ? buffer_6_destinationRegister : _GEN_69; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_71 = 4'h7 == index ? buffer_7_destinationRegister : _GEN_70; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_72 = 4'h8 == index ? buffer_8_destinationRegister : _GEN_71; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_73 = 4'h9 == index ? buffer_9_destinationRegister : _GEN_72; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_74 = 4'ha == index ? buffer_10_destinationRegister : _GEN_73; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_75 = 4'hb == index ? buffer_11_destinationRegister : _GEN_74; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_76 = 4'hc == index ? buffer_12_destinationRegister : _GEN_75; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_77 = 4'hd == index ? buffer_13_destinationRegister : _GEN_76; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_78 = 4'he == index ? buffer_14_destinationRegister : _GEN_77; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_79 = 4'hf == index ? buffer_15_destinationRegister : _GEN_78; // @[ReorderBuffer.scala 91:{37,37}]
  wire [3:0] _GEN_81 = 5'h1 == _GEN_79 ? registerTagMap_1_tagId : 4'h0; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_82 = 5'h2 == _GEN_79 ? registerTagMap_2_tagId : _GEN_81; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_83 = 5'h3 == _GEN_79 ? registerTagMap_3_tagId : _GEN_82; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_84 = 5'h4 == _GEN_79 ? registerTagMap_4_tagId : _GEN_83; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_85 = 5'h5 == _GEN_79 ? registerTagMap_5_tagId : _GEN_84; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_86 = 5'h6 == _GEN_79 ? registerTagMap_6_tagId : _GEN_85; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_87 = 5'h7 == _GEN_79 ? registerTagMap_7_tagId : _GEN_86; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_88 = 5'h8 == _GEN_79 ? registerTagMap_8_tagId : _GEN_87; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_89 = 5'h9 == _GEN_79 ? registerTagMap_9_tagId : _GEN_88; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_90 = 5'ha == _GEN_79 ? registerTagMap_10_tagId : _GEN_89; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_91 = 5'hb == _GEN_79 ? registerTagMap_11_tagId : _GEN_90; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_92 = 5'hc == _GEN_79 ? registerTagMap_12_tagId : _GEN_91; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_93 = 5'hd == _GEN_79 ? registerTagMap_13_tagId : _GEN_92; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_94 = 5'he == _GEN_79 ? registerTagMap_14_tagId : _GEN_93; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_95 = 5'hf == _GEN_79 ? registerTagMap_15_tagId : _GEN_94; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_96 = 5'h10 == _GEN_79 ? registerTagMap_16_tagId : _GEN_95; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_97 = 5'h11 == _GEN_79 ? registerTagMap_17_tagId : _GEN_96; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_98 = 5'h12 == _GEN_79 ? registerTagMap_18_tagId : _GEN_97; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_99 = 5'h13 == _GEN_79 ? registerTagMap_19_tagId : _GEN_98; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_100 = 5'h14 == _GEN_79 ? registerTagMap_20_tagId : _GEN_99; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_101 = 5'h15 == _GEN_79 ? registerTagMap_21_tagId : _GEN_100; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_102 = 5'h16 == _GEN_79 ? registerTagMap_22_tagId : _GEN_101; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_103 = 5'h17 == _GEN_79 ? registerTagMap_23_tagId : _GEN_102; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_104 = 5'h18 == _GEN_79 ? registerTagMap_24_tagId : _GEN_103; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_105 = 5'h19 == _GEN_79 ? registerTagMap_25_tagId : _GEN_104; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_106 = 5'h1a == _GEN_79 ? registerTagMap_26_tagId : _GEN_105; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_107 = 5'h1b == _GEN_79 ? registerTagMap_27_tagId : _GEN_106; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_108 = 5'h1c == _GEN_79 ? registerTagMap_28_tagId : _GEN_107; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_109 = 5'h1d == _GEN_79 ? registerTagMap_29_tagId : _GEN_108; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_110 = 5'h1e == _GEN_79 ? registerTagMap_30_tagId : _GEN_109; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_111 = 5'h1f == _GEN_79 ? registerTagMap_31_tagId : _GEN_110; // @[ReorderBuffer.scala 93:{17,17}]
  wire  _T_1 = index == _GEN_111; // @[ReorderBuffer.scala 93:17]
  wire  _GEN_145 = 5'h1 == _GEN_79 ? 1'h0 : registerTagMap_1_valid; // @[ReorderBuffer.scala 97:{13,13} 69:39]
  wire  _GEN_146 = 5'h2 == _GEN_79 ? 1'h0 : registerTagMap_2_valid; // @[ReorderBuffer.scala 97:{13,13} 69:39]
  wire  _GEN_147 = 5'h3 == _GEN_79 ? 1'h0 : registerTagMap_3_valid; // @[ReorderBuffer.scala 97:{13,13} 69:39]
  wire  _GEN_148 = 5'h4 == _GEN_79 ? 1'h0 : registerTagMap_4_valid; // @[ReorderBuffer.scala 97:{13,13} 69:39]
  wire  _GEN_149 = 5'h5 == _GEN_79 ? 1'h0 : registerTagMap_5_valid; // @[ReorderBuffer.scala 97:{13,13} 69:39]
  wire  _GEN_150 = 5'h6 == _GEN_79 ? 1'h0 : registerTagMap_6_valid; // @[ReorderBuffer.scala 97:{13,13} 69:39]
  wire  _GEN_151 = 5'h7 == _GEN_79 ? 1'h0 : registerTagMap_7_valid; // @[ReorderBuffer.scala 97:{13,13} 69:39]
  wire  _GEN_152 = 5'h8 == _GEN_79 ? 1'h0 : registerTagMap_8_valid; // @[ReorderBuffer.scala 97:{13,13} 69:39]
  wire  _GEN_153 = 5'h9 == _GEN_79 ? 1'h0 : registerTagMap_9_valid; // @[ReorderBuffer.scala 97:{13,13} 69:39]
  wire  _GEN_154 = 5'ha == _GEN_79 ? 1'h0 : registerTagMap_10_valid; // @[ReorderBuffer.scala 97:{13,13} 69:39]
  wire  _GEN_155 = 5'hb == _GEN_79 ? 1'h0 : registerTagMap_11_valid; // @[ReorderBuffer.scala 97:{13,13} 69:39]
  wire  _GEN_156 = 5'hc == _GEN_79 ? 1'h0 : registerTagMap_12_valid; // @[ReorderBuffer.scala 97:{13,13} 69:39]
  wire  _GEN_157 = 5'hd == _GEN_79 ? 1'h0 : registerTagMap_13_valid; // @[ReorderBuffer.scala 97:{13,13} 69:39]
  wire  _GEN_158 = 5'he == _GEN_79 ? 1'h0 : registerTagMap_14_valid; // @[ReorderBuffer.scala 97:{13,13} 69:39]
  wire  _GEN_159 = 5'hf == _GEN_79 ? 1'h0 : registerTagMap_15_valid; // @[ReorderBuffer.scala 97:{13,13} 69:39]
  wire  _GEN_160 = 5'h10 == _GEN_79 ? 1'h0 : registerTagMap_16_valid; // @[ReorderBuffer.scala 97:{13,13} 69:39]
  wire  _GEN_161 = 5'h11 == _GEN_79 ? 1'h0 : registerTagMap_17_valid; // @[ReorderBuffer.scala 97:{13,13} 69:39]
  wire  _GEN_162 = 5'h12 == _GEN_79 ? 1'h0 : registerTagMap_18_valid; // @[ReorderBuffer.scala 97:{13,13} 69:39]
  wire  _GEN_163 = 5'h13 == _GEN_79 ? 1'h0 : registerTagMap_19_valid; // @[ReorderBuffer.scala 97:{13,13} 69:39]
  wire  _GEN_164 = 5'h14 == _GEN_79 ? 1'h0 : registerTagMap_20_valid; // @[ReorderBuffer.scala 97:{13,13} 69:39]
  wire  _GEN_165 = 5'h15 == _GEN_79 ? 1'h0 : registerTagMap_21_valid; // @[ReorderBuffer.scala 97:{13,13} 69:39]
  wire  _GEN_166 = 5'h16 == _GEN_79 ? 1'h0 : registerTagMap_22_valid; // @[ReorderBuffer.scala 97:{13,13} 69:39]
  wire  _GEN_167 = 5'h17 == _GEN_79 ? 1'h0 : registerTagMap_23_valid; // @[ReorderBuffer.scala 97:{13,13} 69:39]
  wire  _GEN_168 = 5'h18 == _GEN_79 ? 1'h0 : registerTagMap_24_valid; // @[ReorderBuffer.scala 97:{13,13} 69:39]
  wire  _GEN_169 = 5'h19 == _GEN_79 ? 1'h0 : registerTagMap_25_valid; // @[ReorderBuffer.scala 97:{13,13} 69:39]
  wire  _GEN_170 = 5'h1a == _GEN_79 ? 1'h0 : registerTagMap_26_valid; // @[ReorderBuffer.scala 97:{13,13} 69:39]
  wire  _GEN_171 = 5'h1b == _GEN_79 ? 1'h0 : registerTagMap_27_valid; // @[ReorderBuffer.scala 97:{13,13} 69:39]
  wire  _GEN_172 = 5'h1c == _GEN_79 ? 1'h0 : registerTagMap_28_valid; // @[ReorderBuffer.scala 97:{13,13} 69:39]
  wire  _GEN_173 = 5'h1d == _GEN_79 ? 1'h0 : registerTagMap_29_valid; // @[ReorderBuffer.scala 97:{13,13} 69:39]
  wire  _GEN_174 = 5'h1e == _GEN_79 ? 1'h0 : registerTagMap_30_valid; // @[ReorderBuffer.scala 97:{13,13} 69:39]
  wire  _GEN_175 = 5'h1f == _GEN_79 ? 1'h0 : registerTagMap_31_valid; // @[ReorderBuffer.scala 97:{13,13} 69:39]
  wire  _GEN_177 = _T_1 ? _GEN_145 : registerTagMap_1_valid; // @[ReorderBuffer.scala 94:11 69:39]
  wire  _GEN_178 = _T_1 ? _GEN_146 : registerTagMap_2_valid; // @[ReorderBuffer.scala 94:11 69:39]
  wire  _GEN_179 = _T_1 ? _GEN_147 : registerTagMap_3_valid; // @[ReorderBuffer.scala 94:11 69:39]
  wire  _GEN_180 = _T_1 ? _GEN_148 : registerTagMap_4_valid; // @[ReorderBuffer.scala 94:11 69:39]
  wire  _GEN_181 = _T_1 ? _GEN_149 : registerTagMap_5_valid; // @[ReorderBuffer.scala 94:11 69:39]
  wire  _GEN_182 = _T_1 ? _GEN_150 : registerTagMap_6_valid; // @[ReorderBuffer.scala 94:11 69:39]
  wire  _GEN_183 = _T_1 ? _GEN_151 : registerTagMap_7_valid; // @[ReorderBuffer.scala 94:11 69:39]
  wire  _GEN_184 = _T_1 ? _GEN_152 : registerTagMap_8_valid; // @[ReorderBuffer.scala 94:11 69:39]
  wire  _GEN_185 = _T_1 ? _GEN_153 : registerTagMap_9_valid; // @[ReorderBuffer.scala 94:11 69:39]
  wire  _GEN_186 = _T_1 ? _GEN_154 : registerTagMap_10_valid; // @[ReorderBuffer.scala 94:11 69:39]
  wire  _GEN_187 = _T_1 ? _GEN_155 : registerTagMap_11_valid; // @[ReorderBuffer.scala 94:11 69:39]
  wire  _GEN_188 = _T_1 ? _GEN_156 : registerTagMap_12_valid; // @[ReorderBuffer.scala 94:11 69:39]
  wire  _GEN_189 = _T_1 ? _GEN_157 : registerTagMap_13_valid; // @[ReorderBuffer.scala 94:11 69:39]
  wire  _GEN_190 = _T_1 ? _GEN_158 : registerTagMap_14_valid; // @[ReorderBuffer.scala 94:11 69:39]
  wire  _GEN_191 = _T_1 ? _GEN_159 : registerTagMap_15_valid; // @[ReorderBuffer.scala 94:11 69:39]
  wire  _GEN_192 = _T_1 ? _GEN_160 : registerTagMap_16_valid; // @[ReorderBuffer.scala 94:11 69:39]
  wire  _GEN_193 = _T_1 ? _GEN_161 : registerTagMap_17_valid; // @[ReorderBuffer.scala 94:11 69:39]
  wire  _GEN_194 = _T_1 ? _GEN_162 : registerTagMap_18_valid; // @[ReorderBuffer.scala 94:11 69:39]
  wire  _GEN_195 = _T_1 ? _GEN_163 : registerTagMap_19_valid; // @[ReorderBuffer.scala 94:11 69:39]
  wire  _GEN_196 = _T_1 ? _GEN_164 : registerTagMap_20_valid; // @[ReorderBuffer.scala 94:11 69:39]
  wire  _GEN_197 = _T_1 ? _GEN_165 : registerTagMap_21_valid; // @[ReorderBuffer.scala 94:11 69:39]
  wire  _GEN_198 = _T_1 ? _GEN_166 : registerTagMap_22_valid; // @[ReorderBuffer.scala 94:11 69:39]
  wire  _GEN_199 = _T_1 ? _GEN_167 : registerTagMap_23_valid; // @[ReorderBuffer.scala 94:11 69:39]
  wire  _GEN_200 = _T_1 ? _GEN_168 : registerTagMap_24_valid; // @[ReorderBuffer.scala 94:11 69:39]
  wire  _GEN_201 = _T_1 ? _GEN_169 : registerTagMap_25_valid; // @[ReorderBuffer.scala 94:11 69:39]
  wire  _GEN_202 = _T_1 ? _GEN_170 : registerTagMap_26_valid; // @[ReorderBuffer.scala 94:11 69:39]
  wire  _GEN_203 = _T_1 ? _GEN_171 : registerTagMap_27_valid; // @[ReorderBuffer.scala 94:11 69:39]
  wire  _GEN_204 = _T_1 ? _GEN_172 : registerTagMap_28_valid; // @[ReorderBuffer.scala 94:11 69:39]
  wire  _GEN_205 = _T_1 ? _GEN_173 : registerTagMap_29_valid; // @[ReorderBuffer.scala 94:11 69:39]
  wire  _GEN_206 = _T_1 ? _GEN_174 : registerTagMap_30_valid; // @[ReorderBuffer.scala 94:11 69:39]
  wire  _GEN_207 = _T_1 ? _GEN_175 : registerTagMap_31_valid; // @[ReorderBuffer.scala 94:11 69:39]
  wire [63:0] _GEN_208 = _io_registerFile_0_valid_T ? _GEN_63 : 64'h0; // @[ReorderBuffer.scala 84:19 89:22 90:23]
  wire [4:0] _GEN_209 = _io_registerFile_0_valid_T ? _GEN_79 : 5'h0; // @[ReorderBuffer.scala 89:22 85:33 91:37]
  wire  _GEN_211 = _io_registerFile_0_valid_T ? _GEN_177 : registerTagMap_1_valid; // @[ReorderBuffer.scala 89:22 69:39]
  wire  _GEN_212 = _io_registerFile_0_valid_T ? _GEN_178 : registerTagMap_2_valid; // @[ReorderBuffer.scala 89:22 69:39]
  wire  _GEN_213 = _io_registerFile_0_valid_T ? _GEN_179 : registerTagMap_3_valid; // @[ReorderBuffer.scala 89:22 69:39]
  wire  _GEN_214 = _io_registerFile_0_valid_T ? _GEN_180 : registerTagMap_4_valid; // @[ReorderBuffer.scala 89:22 69:39]
  wire  _GEN_215 = _io_registerFile_0_valid_T ? _GEN_181 : registerTagMap_5_valid; // @[ReorderBuffer.scala 89:22 69:39]
  wire  _GEN_216 = _io_registerFile_0_valid_T ? _GEN_182 : registerTagMap_6_valid; // @[ReorderBuffer.scala 89:22 69:39]
  wire  _GEN_217 = _io_registerFile_0_valid_T ? _GEN_183 : registerTagMap_7_valid; // @[ReorderBuffer.scala 89:22 69:39]
  wire  _GEN_218 = _io_registerFile_0_valid_T ? _GEN_184 : registerTagMap_8_valid; // @[ReorderBuffer.scala 89:22 69:39]
  wire  _GEN_219 = _io_registerFile_0_valid_T ? _GEN_185 : registerTagMap_9_valid; // @[ReorderBuffer.scala 89:22 69:39]
  wire  _GEN_220 = _io_registerFile_0_valid_T ? _GEN_186 : registerTagMap_10_valid; // @[ReorderBuffer.scala 89:22 69:39]
  wire  _GEN_221 = _io_registerFile_0_valid_T ? _GEN_187 : registerTagMap_11_valid; // @[ReorderBuffer.scala 89:22 69:39]
  wire  _GEN_222 = _io_registerFile_0_valid_T ? _GEN_188 : registerTagMap_12_valid; // @[ReorderBuffer.scala 89:22 69:39]
  wire  _GEN_223 = _io_registerFile_0_valid_T ? _GEN_189 : registerTagMap_13_valid; // @[ReorderBuffer.scala 89:22 69:39]
  wire  _GEN_224 = _io_registerFile_0_valid_T ? _GEN_190 : registerTagMap_14_valid; // @[ReorderBuffer.scala 89:22 69:39]
  wire  _GEN_225 = _io_registerFile_0_valid_T ? _GEN_191 : registerTagMap_15_valid; // @[ReorderBuffer.scala 89:22 69:39]
  wire  _GEN_226 = _io_registerFile_0_valid_T ? _GEN_192 : registerTagMap_16_valid; // @[ReorderBuffer.scala 89:22 69:39]
  wire  _GEN_227 = _io_registerFile_0_valid_T ? _GEN_193 : registerTagMap_17_valid; // @[ReorderBuffer.scala 89:22 69:39]
  wire  _GEN_228 = _io_registerFile_0_valid_T ? _GEN_194 : registerTagMap_18_valid; // @[ReorderBuffer.scala 89:22 69:39]
  wire  _GEN_229 = _io_registerFile_0_valid_T ? _GEN_195 : registerTagMap_19_valid; // @[ReorderBuffer.scala 89:22 69:39]
  wire  _GEN_230 = _io_registerFile_0_valid_T ? _GEN_196 : registerTagMap_20_valid; // @[ReorderBuffer.scala 89:22 69:39]
  wire  _GEN_231 = _io_registerFile_0_valid_T ? _GEN_197 : registerTagMap_21_valid; // @[ReorderBuffer.scala 89:22 69:39]
  wire  _GEN_232 = _io_registerFile_0_valid_T ? _GEN_198 : registerTagMap_22_valid; // @[ReorderBuffer.scala 89:22 69:39]
  wire  _GEN_233 = _io_registerFile_0_valid_T ? _GEN_199 : registerTagMap_23_valid; // @[ReorderBuffer.scala 89:22 69:39]
  wire  _GEN_234 = _io_registerFile_0_valid_T ? _GEN_200 : registerTagMap_24_valid; // @[ReorderBuffer.scala 89:22 69:39]
  wire  _GEN_235 = _io_registerFile_0_valid_T ? _GEN_201 : registerTagMap_25_valid; // @[ReorderBuffer.scala 89:22 69:39]
  wire  _GEN_236 = _io_registerFile_0_valid_T ? _GEN_202 : registerTagMap_26_valid; // @[ReorderBuffer.scala 89:22 69:39]
  wire  _GEN_237 = _io_registerFile_0_valid_T ? _GEN_203 : registerTagMap_27_valid; // @[ReorderBuffer.scala 89:22 69:39]
  wire  _GEN_238 = _io_registerFile_0_valid_T ? _GEN_204 : registerTagMap_28_valid; // @[ReorderBuffer.scala 89:22 69:39]
  wire  _GEN_239 = _io_registerFile_0_valid_T ? _GEN_205 : registerTagMap_29_valid; // @[ReorderBuffer.scala 89:22 69:39]
  wire  _GEN_240 = _io_registerFile_0_valid_T ? _GEN_206 : registerTagMap_30_valid; // @[ReorderBuffer.scala 89:22 69:39]
  wire  _GEN_241 = _io_registerFile_0_valid_T ? _GEN_207 : registerTagMap_31_valid; // @[ReorderBuffer.scala 89:22 69:39]
  wire  _GEN_242 = _io_registerFile_0_valid_T ? 1'h0 : 1'h1; // @[ReorderBuffer.scala 89:22 86:25 100:29]
  wire  _GEN_247 = canCommit ? _GEN_211 : registerTagMap_1_valid; // @[ReorderBuffer.scala 88:21 69:39]
  wire  _GEN_248 = canCommit ? _GEN_212 : registerTagMap_2_valid; // @[ReorderBuffer.scala 88:21 69:39]
  wire  _GEN_249 = canCommit ? _GEN_213 : registerTagMap_3_valid; // @[ReorderBuffer.scala 88:21 69:39]
  wire  _GEN_250 = canCommit ? _GEN_214 : registerTagMap_4_valid; // @[ReorderBuffer.scala 88:21 69:39]
  wire  _GEN_251 = canCommit ? _GEN_215 : registerTagMap_5_valid; // @[ReorderBuffer.scala 88:21 69:39]
  wire  _GEN_252 = canCommit ? _GEN_216 : registerTagMap_6_valid; // @[ReorderBuffer.scala 88:21 69:39]
  wire  _GEN_253 = canCommit ? _GEN_217 : registerTagMap_7_valid; // @[ReorderBuffer.scala 88:21 69:39]
  wire  _GEN_254 = canCommit ? _GEN_218 : registerTagMap_8_valid; // @[ReorderBuffer.scala 88:21 69:39]
  wire  _GEN_255 = canCommit ? _GEN_219 : registerTagMap_9_valid; // @[ReorderBuffer.scala 88:21 69:39]
  wire  _GEN_256 = canCommit ? _GEN_220 : registerTagMap_10_valid; // @[ReorderBuffer.scala 88:21 69:39]
  wire  _GEN_257 = canCommit ? _GEN_221 : registerTagMap_11_valid; // @[ReorderBuffer.scala 88:21 69:39]
  wire  _GEN_258 = canCommit ? _GEN_222 : registerTagMap_12_valid; // @[ReorderBuffer.scala 88:21 69:39]
  wire  _GEN_259 = canCommit ? _GEN_223 : registerTagMap_13_valid; // @[ReorderBuffer.scala 88:21 69:39]
  wire  _GEN_260 = canCommit ? _GEN_224 : registerTagMap_14_valid; // @[ReorderBuffer.scala 88:21 69:39]
  wire  _GEN_261 = canCommit ? _GEN_225 : registerTagMap_15_valid; // @[ReorderBuffer.scala 88:21 69:39]
  wire  _GEN_262 = canCommit ? _GEN_226 : registerTagMap_16_valid; // @[ReorderBuffer.scala 88:21 69:39]
  wire  _GEN_263 = canCommit ? _GEN_227 : registerTagMap_17_valid; // @[ReorderBuffer.scala 88:21 69:39]
  wire  _GEN_264 = canCommit ? _GEN_228 : registerTagMap_18_valid; // @[ReorderBuffer.scala 88:21 69:39]
  wire  _GEN_265 = canCommit ? _GEN_229 : registerTagMap_19_valid; // @[ReorderBuffer.scala 88:21 69:39]
  wire  _GEN_266 = canCommit ? _GEN_230 : registerTagMap_20_valid; // @[ReorderBuffer.scala 88:21 69:39]
  wire  _GEN_267 = canCommit ? _GEN_231 : registerTagMap_21_valid; // @[ReorderBuffer.scala 88:21 69:39]
  wire  _GEN_268 = canCommit ? _GEN_232 : registerTagMap_22_valid; // @[ReorderBuffer.scala 88:21 69:39]
  wire  _GEN_269 = canCommit ? _GEN_233 : registerTagMap_23_valid; // @[ReorderBuffer.scala 88:21 69:39]
  wire  _GEN_270 = canCommit ? _GEN_234 : registerTagMap_24_valid; // @[ReorderBuffer.scala 88:21 69:39]
  wire  _GEN_271 = canCommit ? _GEN_235 : registerTagMap_25_valid; // @[ReorderBuffer.scala 88:21 69:39]
  wire  _GEN_272 = canCommit ? _GEN_236 : registerTagMap_26_valid; // @[ReorderBuffer.scala 88:21 69:39]
  wire  _GEN_273 = canCommit ? _GEN_237 : registerTagMap_27_valid; // @[ReorderBuffer.scala 88:21 69:39]
  wire  _GEN_274 = canCommit ? _GEN_238 : registerTagMap_28_valid; // @[ReorderBuffer.scala 88:21 69:39]
  wire  _GEN_275 = canCommit ? _GEN_239 : registerTagMap_29_valid; // @[ReorderBuffer.scala 88:21 69:39]
  wire  _GEN_276 = canCommit ? _GEN_240 : registerTagMap_30_valid; // @[ReorderBuffer.scala 88:21 69:39]
  wire  _GEN_277 = canCommit ? _GEN_241 : registerTagMap_31_valid; // @[ReorderBuffer.scala 88:21 69:39]
  wire  _GEN_278 = canCommit & _GEN_242; // @[ReorderBuffer.scala 88:21 86:25]
  wire [3:0] index_1 = tail + 4'h1; // @[ReorderBuffer.scala 77:22]
  wire  _GEN_300 = 4'h1 == index_1 ? buffer_1_valueReady : buffer_0_valueReady; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_301 = 4'h2 == index_1 ? buffer_2_valueReady : _GEN_300; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_302 = 4'h3 == index_1 ? buffer_3_valueReady : _GEN_301; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_303 = 4'h4 == index_1 ? buffer_4_valueReady : _GEN_302; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_304 = 4'h5 == index_1 ? buffer_5_valueReady : _GEN_303; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_305 = 4'h6 == index_1 ? buffer_6_valueReady : _GEN_304; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_306 = 4'h7 == index_1 ? buffer_7_valueReady : _GEN_305; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_307 = 4'h8 == index_1 ? buffer_8_valueReady : _GEN_306; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_308 = 4'h9 == index_1 ? buffer_9_valueReady : _GEN_307; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_309 = 4'ha == index_1 ? buffer_10_valueReady : _GEN_308; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_310 = 4'hb == index_1 ? buffer_11_valueReady : _GEN_309; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_311 = 4'hc == index_1 ? buffer_12_valueReady : _GEN_310; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_312 = 4'hd == index_1 ? buffer_13_valueReady : _GEN_311; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_313 = 4'he == index_1 ? buffer_14_valueReady : _GEN_312; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_314 = 4'hf == index_1 ? buffer_15_valueReady : _GEN_313; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_316 = 4'h1 == index_1 ? buffer_1_storeSign : buffer_0_storeSign; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_317 = 4'h2 == index_1 ? buffer_2_storeSign : _GEN_316; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_318 = 4'h3 == index_1 ? buffer_3_storeSign : _GEN_317; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_319 = 4'h4 == index_1 ? buffer_4_storeSign : _GEN_318; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_320 = 4'h5 == index_1 ? buffer_5_storeSign : _GEN_319; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_321 = 4'h6 == index_1 ? buffer_6_storeSign : _GEN_320; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_322 = 4'h7 == index_1 ? buffer_7_storeSign : _GEN_321; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_323 = 4'h8 == index_1 ? buffer_8_storeSign : _GEN_322; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_324 = 4'h9 == index_1 ? buffer_9_storeSign : _GEN_323; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_325 = 4'ha == index_1 ? buffer_10_storeSign : _GEN_324; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_326 = 4'hb == index_1 ? buffer_11_storeSign : _GEN_325; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_327 = 4'hc == index_1 ? buffer_12_storeSign : _GEN_326; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_328 = 4'hd == index_1 ? buffer_13_storeSign : _GEN_327; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_329 = 4'he == index_1 ? buffer_14_storeSign : _GEN_328; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_330 = 4'hf == index_1 ? buffer_15_storeSign : _GEN_329; // @[ReorderBuffer.scala 79:{50,50}]
  wire  instructionOk_1 = _GEN_314 | _GEN_330; // @[ReorderBuffer.scala 79:50]
  wire  canCommit_1 = canCommit & index_1 != head & instructionOk_1; // @[ReorderBuffer.scala 80:49]
  wire  _GEN_332 = 4'h1 == index_1 ? buffer_1_isError : buffer_0_isError; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_333 = 4'h2 == index_1 ? buffer_2_isError : _GEN_332; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_334 = 4'h3 == index_1 ? buffer_3_isError : _GEN_333; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_335 = 4'h4 == index_1 ? buffer_4_isError : _GEN_334; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_336 = 4'h5 == index_1 ? buffer_5_isError : _GEN_335; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_337 = 4'h6 == index_1 ? buffer_6_isError : _GEN_336; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_338 = 4'h7 == index_1 ? buffer_7_isError : _GEN_337; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_339 = 4'h8 == index_1 ? buffer_8_isError : _GEN_338; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_340 = 4'h9 == index_1 ? buffer_9_isError : _GEN_339; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_341 = 4'ha == index_1 ? buffer_10_isError : _GEN_340; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_342 = 4'hb == index_1 ? buffer_11_isError : _GEN_341; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_343 = 4'hc == index_1 ? buffer_12_isError : _GEN_342; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_344 = 4'hd == index_1 ? buffer_13_isError : _GEN_343; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_345 = 4'he == index_1 ? buffer_14_isError : _GEN_344; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_346 = 4'hf == index_1 ? buffer_15_isError : _GEN_345; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _io_registerFile_1_valid_T = ~_GEN_346; // @[ReorderBuffer.scala 83:30]
  wire [63:0] _GEN_348 = 4'h1 == index_1 ? buffer_1_value : buffer_0_value; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_349 = 4'h2 == index_1 ? buffer_2_value : _GEN_348; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_350 = 4'h3 == index_1 ? buffer_3_value : _GEN_349; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_351 = 4'h4 == index_1 ? buffer_4_value : _GEN_350; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_352 = 4'h5 == index_1 ? buffer_5_value : _GEN_351; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_353 = 4'h6 == index_1 ? buffer_6_value : _GEN_352; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_354 = 4'h7 == index_1 ? buffer_7_value : _GEN_353; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_355 = 4'h8 == index_1 ? buffer_8_value : _GEN_354; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_356 = 4'h9 == index_1 ? buffer_9_value : _GEN_355; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_357 = 4'ha == index_1 ? buffer_10_value : _GEN_356; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_358 = 4'hb == index_1 ? buffer_11_value : _GEN_357; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_359 = 4'hc == index_1 ? buffer_12_value : _GEN_358; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_360 = 4'hd == index_1 ? buffer_13_value : _GEN_359; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_361 = 4'he == index_1 ? buffer_14_value : _GEN_360; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_362 = 4'hf == index_1 ? buffer_15_value : _GEN_361; // @[ReorderBuffer.scala 90:{23,23}]
  wire [4:0] _GEN_364 = 4'h1 == index_1 ? buffer_1_destinationRegister : buffer_0_destinationRegister; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_365 = 4'h2 == index_1 ? buffer_2_destinationRegister : _GEN_364; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_366 = 4'h3 == index_1 ? buffer_3_destinationRegister : _GEN_365; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_367 = 4'h4 == index_1 ? buffer_4_destinationRegister : _GEN_366; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_368 = 4'h5 == index_1 ? buffer_5_destinationRegister : _GEN_367; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_369 = 4'h6 == index_1 ? buffer_6_destinationRegister : _GEN_368; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_370 = 4'h7 == index_1 ? buffer_7_destinationRegister : _GEN_369; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_371 = 4'h8 == index_1 ? buffer_8_destinationRegister : _GEN_370; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_372 = 4'h9 == index_1 ? buffer_9_destinationRegister : _GEN_371; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_373 = 4'ha == index_1 ? buffer_10_destinationRegister : _GEN_372; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_374 = 4'hb == index_1 ? buffer_11_destinationRegister : _GEN_373; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_375 = 4'hc == index_1 ? buffer_12_destinationRegister : _GEN_374; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_376 = 4'hd == index_1 ? buffer_13_destinationRegister : _GEN_375; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_377 = 4'he == index_1 ? buffer_14_destinationRegister : _GEN_376; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_378 = 4'hf == index_1 ? buffer_15_destinationRegister : _GEN_377; // @[ReorderBuffer.scala 91:{37,37}]
  wire [3:0] _GEN_380 = 5'h1 == _GEN_378 ? registerTagMap_1_tagId : 4'h0; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_381 = 5'h2 == _GEN_378 ? registerTagMap_2_tagId : _GEN_380; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_382 = 5'h3 == _GEN_378 ? registerTagMap_3_tagId : _GEN_381; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_383 = 5'h4 == _GEN_378 ? registerTagMap_4_tagId : _GEN_382; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_384 = 5'h5 == _GEN_378 ? registerTagMap_5_tagId : _GEN_383; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_385 = 5'h6 == _GEN_378 ? registerTagMap_6_tagId : _GEN_384; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_386 = 5'h7 == _GEN_378 ? registerTagMap_7_tagId : _GEN_385; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_387 = 5'h8 == _GEN_378 ? registerTagMap_8_tagId : _GEN_386; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_388 = 5'h9 == _GEN_378 ? registerTagMap_9_tagId : _GEN_387; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_389 = 5'ha == _GEN_378 ? registerTagMap_10_tagId : _GEN_388; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_390 = 5'hb == _GEN_378 ? registerTagMap_11_tagId : _GEN_389; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_391 = 5'hc == _GEN_378 ? registerTagMap_12_tagId : _GEN_390; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_392 = 5'hd == _GEN_378 ? registerTagMap_13_tagId : _GEN_391; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_393 = 5'he == _GEN_378 ? registerTagMap_14_tagId : _GEN_392; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_394 = 5'hf == _GEN_378 ? registerTagMap_15_tagId : _GEN_393; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_395 = 5'h10 == _GEN_378 ? registerTagMap_16_tagId : _GEN_394; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_396 = 5'h11 == _GEN_378 ? registerTagMap_17_tagId : _GEN_395; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_397 = 5'h12 == _GEN_378 ? registerTagMap_18_tagId : _GEN_396; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_398 = 5'h13 == _GEN_378 ? registerTagMap_19_tagId : _GEN_397; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_399 = 5'h14 == _GEN_378 ? registerTagMap_20_tagId : _GEN_398; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_400 = 5'h15 == _GEN_378 ? registerTagMap_21_tagId : _GEN_399; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_401 = 5'h16 == _GEN_378 ? registerTagMap_22_tagId : _GEN_400; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_402 = 5'h17 == _GEN_378 ? registerTagMap_23_tagId : _GEN_401; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_403 = 5'h18 == _GEN_378 ? registerTagMap_24_tagId : _GEN_402; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_404 = 5'h19 == _GEN_378 ? registerTagMap_25_tagId : _GEN_403; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_405 = 5'h1a == _GEN_378 ? registerTagMap_26_tagId : _GEN_404; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_406 = 5'h1b == _GEN_378 ? registerTagMap_27_tagId : _GEN_405; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_407 = 5'h1c == _GEN_378 ? registerTagMap_28_tagId : _GEN_406; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_408 = 5'h1d == _GEN_378 ? registerTagMap_29_tagId : _GEN_407; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_409 = 5'h1e == _GEN_378 ? registerTagMap_30_tagId : _GEN_408; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_410 = 5'h1f == _GEN_378 ? registerTagMap_31_tagId : _GEN_409; // @[ReorderBuffer.scala 93:{17,17}]
  wire  _T_3 = index_1 == _GEN_410; // @[ReorderBuffer.scala 93:17]
  wire  _GEN_444 = 5'h1 == _GEN_378 ? 1'h0 : _GEN_247; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_445 = 5'h2 == _GEN_378 ? 1'h0 : _GEN_248; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_446 = 5'h3 == _GEN_378 ? 1'h0 : _GEN_249; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_447 = 5'h4 == _GEN_378 ? 1'h0 : _GEN_250; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_448 = 5'h5 == _GEN_378 ? 1'h0 : _GEN_251; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_449 = 5'h6 == _GEN_378 ? 1'h0 : _GEN_252; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_450 = 5'h7 == _GEN_378 ? 1'h0 : _GEN_253; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_451 = 5'h8 == _GEN_378 ? 1'h0 : _GEN_254; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_452 = 5'h9 == _GEN_378 ? 1'h0 : _GEN_255; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_453 = 5'ha == _GEN_378 ? 1'h0 : _GEN_256; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_454 = 5'hb == _GEN_378 ? 1'h0 : _GEN_257; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_455 = 5'hc == _GEN_378 ? 1'h0 : _GEN_258; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_456 = 5'hd == _GEN_378 ? 1'h0 : _GEN_259; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_457 = 5'he == _GEN_378 ? 1'h0 : _GEN_260; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_458 = 5'hf == _GEN_378 ? 1'h0 : _GEN_261; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_459 = 5'h10 == _GEN_378 ? 1'h0 : _GEN_262; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_460 = 5'h11 == _GEN_378 ? 1'h0 : _GEN_263; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_461 = 5'h12 == _GEN_378 ? 1'h0 : _GEN_264; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_462 = 5'h13 == _GEN_378 ? 1'h0 : _GEN_265; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_463 = 5'h14 == _GEN_378 ? 1'h0 : _GEN_266; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_464 = 5'h15 == _GEN_378 ? 1'h0 : _GEN_267; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_465 = 5'h16 == _GEN_378 ? 1'h0 : _GEN_268; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_466 = 5'h17 == _GEN_378 ? 1'h0 : _GEN_269; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_467 = 5'h18 == _GEN_378 ? 1'h0 : _GEN_270; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_468 = 5'h19 == _GEN_378 ? 1'h0 : _GEN_271; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_469 = 5'h1a == _GEN_378 ? 1'h0 : _GEN_272; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_470 = 5'h1b == _GEN_378 ? 1'h0 : _GEN_273; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_471 = 5'h1c == _GEN_378 ? 1'h0 : _GEN_274; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_472 = 5'h1d == _GEN_378 ? 1'h0 : _GEN_275; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_473 = 5'h1e == _GEN_378 ? 1'h0 : _GEN_276; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_474 = 5'h1f == _GEN_378 ? 1'h0 : _GEN_277; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_476 = _T_3 ? _GEN_444 : _GEN_247; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_477 = _T_3 ? _GEN_445 : _GEN_248; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_478 = _T_3 ? _GEN_446 : _GEN_249; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_479 = _T_3 ? _GEN_447 : _GEN_250; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_480 = _T_3 ? _GEN_448 : _GEN_251; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_481 = _T_3 ? _GEN_449 : _GEN_252; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_482 = _T_3 ? _GEN_450 : _GEN_253; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_483 = _T_3 ? _GEN_451 : _GEN_254; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_484 = _T_3 ? _GEN_452 : _GEN_255; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_485 = _T_3 ? _GEN_453 : _GEN_256; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_486 = _T_3 ? _GEN_454 : _GEN_257; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_487 = _T_3 ? _GEN_455 : _GEN_258; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_488 = _T_3 ? _GEN_456 : _GEN_259; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_489 = _T_3 ? _GEN_457 : _GEN_260; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_490 = _T_3 ? _GEN_458 : _GEN_261; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_491 = _T_3 ? _GEN_459 : _GEN_262; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_492 = _T_3 ? _GEN_460 : _GEN_263; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_493 = _T_3 ? _GEN_461 : _GEN_264; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_494 = _T_3 ? _GEN_462 : _GEN_265; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_495 = _T_3 ? _GEN_463 : _GEN_266; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_496 = _T_3 ? _GEN_464 : _GEN_267; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_497 = _T_3 ? _GEN_465 : _GEN_268; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_498 = _T_3 ? _GEN_466 : _GEN_269; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_499 = _T_3 ? _GEN_467 : _GEN_270; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_500 = _T_3 ? _GEN_468 : _GEN_271; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_501 = _T_3 ? _GEN_469 : _GEN_272; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_502 = _T_3 ? _GEN_470 : _GEN_273; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_503 = _T_3 ? _GEN_471 : _GEN_274; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_504 = _T_3 ? _GEN_472 : _GEN_275; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_505 = _T_3 ? _GEN_473 : _GEN_276; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_506 = _T_3 ? _GEN_474 : _GEN_277; // @[ReorderBuffer.scala 94:11]
  wire [63:0] _GEN_507 = _io_registerFile_1_valid_T ? _GEN_362 : 64'h0; // @[ReorderBuffer.scala 84:19 89:22 90:23]
  wire [4:0] _GEN_508 = _io_registerFile_1_valid_T ? _GEN_378 : 5'h0; // @[ReorderBuffer.scala 89:22 85:33 91:37]
  wire  _GEN_510 = _io_registerFile_1_valid_T ? _GEN_476 : _GEN_247; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_511 = _io_registerFile_1_valid_T ? _GEN_477 : _GEN_248; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_512 = _io_registerFile_1_valid_T ? _GEN_478 : _GEN_249; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_513 = _io_registerFile_1_valid_T ? _GEN_479 : _GEN_250; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_514 = _io_registerFile_1_valid_T ? _GEN_480 : _GEN_251; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_515 = _io_registerFile_1_valid_T ? _GEN_481 : _GEN_252; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_516 = _io_registerFile_1_valid_T ? _GEN_482 : _GEN_253; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_517 = _io_registerFile_1_valid_T ? _GEN_483 : _GEN_254; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_518 = _io_registerFile_1_valid_T ? _GEN_484 : _GEN_255; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_519 = _io_registerFile_1_valid_T ? _GEN_485 : _GEN_256; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_520 = _io_registerFile_1_valid_T ? _GEN_486 : _GEN_257; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_521 = _io_registerFile_1_valid_T ? _GEN_487 : _GEN_258; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_522 = _io_registerFile_1_valid_T ? _GEN_488 : _GEN_259; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_523 = _io_registerFile_1_valid_T ? _GEN_489 : _GEN_260; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_524 = _io_registerFile_1_valid_T ? _GEN_490 : _GEN_261; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_525 = _io_registerFile_1_valid_T ? _GEN_491 : _GEN_262; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_526 = _io_registerFile_1_valid_T ? _GEN_492 : _GEN_263; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_527 = _io_registerFile_1_valid_T ? _GEN_493 : _GEN_264; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_528 = _io_registerFile_1_valid_T ? _GEN_494 : _GEN_265; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_529 = _io_registerFile_1_valid_T ? _GEN_495 : _GEN_266; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_530 = _io_registerFile_1_valid_T ? _GEN_496 : _GEN_267; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_531 = _io_registerFile_1_valid_T ? _GEN_497 : _GEN_268; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_532 = _io_registerFile_1_valid_T ? _GEN_498 : _GEN_269; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_533 = _io_registerFile_1_valid_T ? _GEN_499 : _GEN_270; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_534 = _io_registerFile_1_valid_T ? _GEN_500 : _GEN_271; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_535 = _io_registerFile_1_valid_T ? _GEN_501 : _GEN_272; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_536 = _io_registerFile_1_valid_T ? _GEN_502 : _GEN_273; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_537 = _io_registerFile_1_valid_T ? _GEN_503 : _GEN_274; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_538 = _io_registerFile_1_valid_T ? _GEN_504 : _GEN_275; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_539 = _io_registerFile_1_valid_T ? _GEN_505 : _GEN_276; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_540 = _io_registerFile_1_valid_T ? _GEN_506 : _GEN_277; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_543 = _io_registerFile_1_valid_T ? _GEN_278 : 1'h1; // @[ReorderBuffer.scala 102:20 89:22]
  wire  _GEN_547 = canCommit_1 ? _GEN_510 : _GEN_247; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_548 = canCommit_1 ? _GEN_511 : _GEN_248; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_549 = canCommit_1 ? _GEN_512 : _GEN_249; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_550 = canCommit_1 ? _GEN_513 : _GEN_250; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_551 = canCommit_1 ? _GEN_514 : _GEN_251; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_552 = canCommit_1 ? _GEN_515 : _GEN_252; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_553 = canCommit_1 ? _GEN_516 : _GEN_253; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_554 = canCommit_1 ? _GEN_517 : _GEN_254; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_555 = canCommit_1 ? _GEN_518 : _GEN_255; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_556 = canCommit_1 ? _GEN_519 : _GEN_256; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_557 = canCommit_1 ? _GEN_520 : _GEN_257; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_558 = canCommit_1 ? _GEN_521 : _GEN_258; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_559 = canCommit_1 ? _GEN_522 : _GEN_259; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_560 = canCommit_1 ? _GEN_523 : _GEN_260; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_561 = canCommit_1 ? _GEN_524 : _GEN_261; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_562 = canCommit_1 ? _GEN_525 : _GEN_262; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_563 = canCommit_1 ? _GEN_526 : _GEN_263; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_564 = canCommit_1 ? _GEN_527 : _GEN_264; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_565 = canCommit_1 ? _GEN_528 : _GEN_265; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_566 = canCommit_1 ? _GEN_529 : _GEN_266; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_567 = canCommit_1 ? _GEN_530 : _GEN_267; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_568 = canCommit_1 ? _GEN_531 : _GEN_268; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_569 = canCommit_1 ? _GEN_532 : _GEN_269; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_570 = canCommit_1 ? _GEN_533 : _GEN_270; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_571 = canCommit_1 ? _GEN_534 : _GEN_271; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_572 = canCommit_1 ? _GEN_535 : _GEN_272; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_573 = canCommit_1 ? _GEN_536 : _GEN_273; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_574 = canCommit_1 ? _GEN_537 : _GEN_274; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_575 = canCommit_1 ? _GEN_538 : _GEN_275; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_576 = canCommit_1 ? _GEN_539 : _GEN_276; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_577 = canCommit_1 ? _GEN_540 : _GEN_277; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_580 = canCommit_1 ? _GEN_543 : _GEN_278; // @[ReorderBuffer.scala 88:21]
  wire [3:0] index_2 = tail + 4'h2; // @[ReorderBuffer.scala 77:22]
  wire  _GEN_601 = 4'h1 == index_2 ? buffer_1_valueReady : buffer_0_valueReady; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_602 = 4'h2 == index_2 ? buffer_2_valueReady : _GEN_601; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_603 = 4'h3 == index_2 ? buffer_3_valueReady : _GEN_602; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_604 = 4'h4 == index_2 ? buffer_4_valueReady : _GEN_603; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_605 = 4'h5 == index_2 ? buffer_5_valueReady : _GEN_604; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_606 = 4'h6 == index_2 ? buffer_6_valueReady : _GEN_605; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_607 = 4'h7 == index_2 ? buffer_7_valueReady : _GEN_606; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_608 = 4'h8 == index_2 ? buffer_8_valueReady : _GEN_607; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_609 = 4'h9 == index_2 ? buffer_9_valueReady : _GEN_608; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_610 = 4'ha == index_2 ? buffer_10_valueReady : _GEN_609; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_611 = 4'hb == index_2 ? buffer_11_valueReady : _GEN_610; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_612 = 4'hc == index_2 ? buffer_12_valueReady : _GEN_611; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_613 = 4'hd == index_2 ? buffer_13_valueReady : _GEN_612; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_614 = 4'he == index_2 ? buffer_14_valueReady : _GEN_613; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_615 = 4'hf == index_2 ? buffer_15_valueReady : _GEN_614; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_617 = 4'h1 == index_2 ? buffer_1_storeSign : buffer_0_storeSign; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_618 = 4'h2 == index_2 ? buffer_2_storeSign : _GEN_617; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_619 = 4'h3 == index_2 ? buffer_3_storeSign : _GEN_618; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_620 = 4'h4 == index_2 ? buffer_4_storeSign : _GEN_619; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_621 = 4'h5 == index_2 ? buffer_5_storeSign : _GEN_620; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_622 = 4'h6 == index_2 ? buffer_6_storeSign : _GEN_621; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_623 = 4'h7 == index_2 ? buffer_7_storeSign : _GEN_622; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_624 = 4'h8 == index_2 ? buffer_8_storeSign : _GEN_623; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_625 = 4'h9 == index_2 ? buffer_9_storeSign : _GEN_624; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_626 = 4'ha == index_2 ? buffer_10_storeSign : _GEN_625; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_627 = 4'hb == index_2 ? buffer_11_storeSign : _GEN_626; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_628 = 4'hc == index_2 ? buffer_12_storeSign : _GEN_627; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_629 = 4'hd == index_2 ? buffer_13_storeSign : _GEN_628; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_630 = 4'he == index_2 ? buffer_14_storeSign : _GEN_629; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_631 = 4'hf == index_2 ? buffer_15_storeSign : _GEN_630; // @[ReorderBuffer.scala 79:{50,50}]
  wire  instructionOk_2 = _GEN_615 | _GEN_631; // @[ReorderBuffer.scala 79:50]
  wire  canCommit_2 = canCommit_1 & index_2 != head & instructionOk_2; // @[ReorderBuffer.scala 80:49]
  wire  _GEN_633 = 4'h1 == index_2 ? buffer_1_isError : buffer_0_isError; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_634 = 4'h2 == index_2 ? buffer_2_isError : _GEN_633; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_635 = 4'h3 == index_2 ? buffer_3_isError : _GEN_634; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_636 = 4'h4 == index_2 ? buffer_4_isError : _GEN_635; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_637 = 4'h5 == index_2 ? buffer_5_isError : _GEN_636; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_638 = 4'h6 == index_2 ? buffer_6_isError : _GEN_637; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_639 = 4'h7 == index_2 ? buffer_7_isError : _GEN_638; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_640 = 4'h8 == index_2 ? buffer_8_isError : _GEN_639; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_641 = 4'h9 == index_2 ? buffer_9_isError : _GEN_640; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_642 = 4'ha == index_2 ? buffer_10_isError : _GEN_641; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_643 = 4'hb == index_2 ? buffer_11_isError : _GEN_642; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_644 = 4'hc == index_2 ? buffer_12_isError : _GEN_643; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_645 = 4'hd == index_2 ? buffer_13_isError : _GEN_644; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_646 = 4'he == index_2 ? buffer_14_isError : _GEN_645; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_647 = 4'hf == index_2 ? buffer_15_isError : _GEN_646; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _io_registerFile_2_valid_T = ~_GEN_647; // @[ReorderBuffer.scala 83:30]
  wire [63:0] _GEN_649 = 4'h1 == index_2 ? buffer_1_value : buffer_0_value; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_650 = 4'h2 == index_2 ? buffer_2_value : _GEN_649; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_651 = 4'h3 == index_2 ? buffer_3_value : _GEN_650; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_652 = 4'h4 == index_2 ? buffer_4_value : _GEN_651; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_653 = 4'h5 == index_2 ? buffer_5_value : _GEN_652; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_654 = 4'h6 == index_2 ? buffer_6_value : _GEN_653; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_655 = 4'h7 == index_2 ? buffer_7_value : _GEN_654; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_656 = 4'h8 == index_2 ? buffer_8_value : _GEN_655; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_657 = 4'h9 == index_2 ? buffer_9_value : _GEN_656; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_658 = 4'ha == index_2 ? buffer_10_value : _GEN_657; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_659 = 4'hb == index_2 ? buffer_11_value : _GEN_658; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_660 = 4'hc == index_2 ? buffer_12_value : _GEN_659; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_661 = 4'hd == index_2 ? buffer_13_value : _GEN_660; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_662 = 4'he == index_2 ? buffer_14_value : _GEN_661; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_663 = 4'hf == index_2 ? buffer_15_value : _GEN_662; // @[ReorderBuffer.scala 90:{23,23}]
  wire [4:0] _GEN_665 = 4'h1 == index_2 ? buffer_1_destinationRegister : buffer_0_destinationRegister; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_666 = 4'h2 == index_2 ? buffer_2_destinationRegister : _GEN_665; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_667 = 4'h3 == index_2 ? buffer_3_destinationRegister : _GEN_666; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_668 = 4'h4 == index_2 ? buffer_4_destinationRegister : _GEN_667; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_669 = 4'h5 == index_2 ? buffer_5_destinationRegister : _GEN_668; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_670 = 4'h6 == index_2 ? buffer_6_destinationRegister : _GEN_669; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_671 = 4'h7 == index_2 ? buffer_7_destinationRegister : _GEN_670; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_672 = 4'h8 == index_2 ? buffer_8_destinationRegister : _GEN_671; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_673 = 4'h9 == index_2 ? buffer_9_destinationRegister : _GEN_672; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_674 = 4'ha == index_2 ? buffer_10_destinationRegister : _GEN_673; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_675 = 4'hb == index_2 ? buffer_11_destinationRegister : _GEN_674; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_676 = 4'hc == index_2 ? buffer_12_destinationRegister : _GEN_675; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_677 = 4'hd == index_2 ? buffer_13_destinationRegister : _GEN_676; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_678 = 4'he == index_2 ? buffer_14_destinationRegister : _GEN_677; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_679 = 4'hf == index_2 ? buffer_15_destinationRegister : _GEN_678; // @[ReorderBuffer.scala 91:{37,37}]
  wire [3:0] _GEN_681 = 5'h1 == _GEN_679 ? registerTagMap_1_tagId : 4'h0; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_682 = 5'h2 == _GEN_679 ? registerTagMap_2_tagId : _GEN_681; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_683 = 5'h3 == _GEN_679 ? registerTagMap_3_tagId : _GEN_682; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_684 = 5'h4 == _GEN_679 ? registerTagMap_4_tagId : _GEN_683; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_685 = 5'h5 == _GEN_679 ? registerTagMap_5_tagId : _GEN_684; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_686 = 5'h6 == _GEN_679 ? registerTagMap_6_tagId : _GEN_685; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_687 = 5'h7 == _GEN_679 ? registerTagMap_7_tagId : _GEN_686; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_688 = 5'h8 == _GEN_679 ? registerTagMap_8_tagId : _GEN_687; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_689 = 5'h9 == _GEN_679 ? registerTagMap_9_tagId : _GEN_688; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_690 = 5'ha == _GEN_679 ? registerTagMap_10_tagId : _GEN_689; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_691 = 5'hb == _GEN_679 ? registerTagMap_11_tagId : _GEN_690; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_692 = 5'hc == _GEN_679 ? registerTagMap_12_tagId : _GEN_691; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_693 = 5'hd == _GEN_679 ? registerTagMap_13_tagId : _GEN_692; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_694 = 5'he == _GEN_679 ? registerTagMap_14_tagId : _GEN_693; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_695 = 5'hf == _GEN_679 ? registerTagMap_15_tagId : _GEN_694; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_696 = 5'h10 == _GEN_679 ? registerTagMap_16_tagId : _GEN_695; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_697 = 5'h11 == _GEN_679 ? registerTagMap_17_tagId : _GEN_696; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_698 = 5'h12 == _GEN_679 ? registerTagMap_18_tagId : _GEN_697; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_699 = 5'h13 == _GEN_679 ? registerTagMap_19_tagId : _GEN_698; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_700 = 5'h14 == _GEN_679 ? registerTagMap_20_tagId : _GEN_699; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_701 = 5'h15 == _GEN_679 ? registerTagMap_21_tagId : _GEN_700; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_702 = 5'h16 == _GEN_679 ? registerTagMap_22_tagId : _GEN_701; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_703 = 5'h17 == _GEN_679 ? registerTagMap_23_tagId : _GEN_702; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_704 = 5'h18 == _GEN_679 ? registerTagMap_24_tagId : _GEN_703; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_705 = 5'h19 == _GEN_679 ? registerTagMap_25_tagId : _GEN_704; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_706 = 5'h1a == _GEN_679 ? registerTagMap_26_tagId : _GEN_705; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_707 = 5'h1b == _GEN_679 ? registerTagMap_27_tagId : _GEN_706; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_708 = 5'h1c == _GEN_679 ? registerTagMap_28_tagId : _GEN_707; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_709 = 5'h1d == _GEN_679 ? registerTagMap_29_tagId : _GEN_708; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_710 = 5'h1e == _GEN_679 ? registerTagMap_30_tagId : _GEN_709; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_711 = 5'h1f == _GEN_679 ? registerTagMap_31_tagId : _GEN_710; // @[ReorderBuffer.scala 93:{17,17}]
  wire  _T_5 = index_2 == _GEN_711; // @[ReorderBuffer.scala 93:17]
  wire  _GEN_745 = 5'h1 == _GEN_679 ? 1'h0 : _GEN_547; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_746 = 5'h2 == _GEN_679 ? 1'h0 : _GEN_548; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_747 = 5'h3 == _GEN_679 ? 1'h0 : _GEN_549; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_748 = 5'h4 == _GEN_679 ? 1'h0 : _GEN_550; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_749 = 5'h5 == _GEN_679 ? 1'h0 : _GEN_551; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_750 = 5'h6 == _GEN_679 ? 1'h0 : _GEN_552; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_751 = 5'h7 == _GEN_679 ? 1'h0 : _GEN_553; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_752 = 5'h8 == _GEN_679 ? 1'h0 : _GEN_554; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_753 = 5'h9 == _GEN_679 ? 1'h0 : _GEN_555; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_754 = 5'ha == _GEN_679 ? 1'h0 : _GEN_556; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_755 = 5'hb == _GEN_679 ? 1'h0 : _GEN_557; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_756 = 5'hc == _GEN_679 ? 1'h0 : _GEN_558; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_757 = 5'hd == _GEN_679 ? 1'h0 : _GEN_559; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_758 = 5'he == _GEN_679 ? 1'h0 : _GEN_560; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_759 = 5'hf == _GEN_679 ? 1'h0 : _GEN_561; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_760 = 5'h10 == _GEN_679 ? 1'h0 : _GEN_562; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_761 = 5'h11 == _GEN_679 ? 1'h0 : _GEN_563; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_762 = 5'h12 == _GEN_679 ? 1'h0 : _GEN_564; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_763 = 5'h13 == _GEN_679 ? 1'h0 : _GEN_565; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_764 = 5'h14 == _GEN_679 ? 1'h0 : _GEN_566; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_765 = 5'h15 == _GEN_679 ? 1'h0 : _GEN_567; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_766 = 5'h16 == _GEN_679 ? 1'h0 : _GEN_568; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_767 = 5'h17 == _GEN_679 ? 1'h0 : _GEN_569; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_768 = 5'h18 == _GEN_679 ? 1'h0 : _GEN_570; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_769 = 5'h19 == _GEN_679 ? 1'h0 : _GEN_571; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_770 = 5'h1a == _GEN_679 ? 1'h0 : _GEN_572; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_771 = 5'h1b == _GEN_679 ? 1'h0 : _GEN_573; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_772 = 5'h1c == _GEN_679 ? 1'h0 : _GEN_574; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_773 = 5'h1d == _GEN_679 ? 1'h0 : _GEN_575; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_774 = 5'h1e == _GEN_679 ? 1'h0 : _GEN_576; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_775 = 5'h1f == _GEN_679 ? 1'h0 : _GEN_577; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_777 = _T_5 ? _GEN_745 : _GEN_547; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_778 = _T_5 ? _GEN_746 : _GEN_548; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_779 = _T_5 ? _GEN_747 : _GEN_549; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_780 = _T_5 ? _GEN_748 : _GEN_550; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_781 = _T_5 ? _GEN_749 : _GEN_551; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_782 = _T_5 ? _GEN_750 : _GEN_552; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_783 = _T_5 ? _GEN_751 : _GEN_553; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_784 = _T_5 ? _GEN_752 : _GEN_554; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_785 = _T_5 ? _GEN_753 : _GEN_555; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_786 = _T_5 ? _GEN_754 : _GEN_556; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_787 = _T_5 ? _GEN_755 : _GEN_557; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_788 = _T_5 ? _GEN_756 : _GEN_558; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_789 = _T_5 ? _GEN_757 : _GEN_559; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_790 = _T_5 ? _GEN_758 : _GEN_560; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_791 = _T_5 ? _GEN_759 : _GEN_561; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_792 = _T_5 ? _GEN_760 : _GEN_562; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_793 = _T_5 ? _GEN_761 : _GEN_563; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_794 = _T_5 ? _GEN_762 : _GEN_564; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_795 = _T_5 ? _GEN_763 : _GEN_565; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_796 = _T_5 ? _GEN_764 : _GEN_566; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_797 = _T_5 ? _GEN_765 : _GEN_567; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_798 = _T_5 ? _GEN_766 : _GEN_568; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_799 = _T_5 ? _GEN_767 : _GEN_569; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_800 = _T_5 ? _GEN_768 : _GEN_570; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_801 = _T_5 ? _GEN_769 : _GEN_571; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_802 = _T_5 ? _GEN_770 : _GEN_572; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_803 = _T_5 ? _GEN_771 : _GEN_573; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_804 = _T_5 ? _GEN_772 : _GEN_574; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_805 = _T_5 ? _GEN_773 : _GEN_575; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_806 = _T_5 ? _GEN_774 : _GEN_576; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_807 = _T_5 ? _GEN_775 : _GEN_577; // @[ReorderBuffer.scala 94:11]
  wire [63:0] _GEN_808 = _io_registerFile_2_valid_T ? _GEN_663 : 64'h0; // @[ReorderBuffer.scala 84:19 89:22 90:23]
  wire [4:0] _GEN_809 = _io_registerFile_2_valid_T ? _GEN_679 : 5'h0; // @[ReorderBuffer.scala 89:22 85:33 91:37]
  wire  _GEN_811 = _io_registerFile_2_valid_T ? _GEN_777 : _GEN_547; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_812 = _io_registerFile_2_valid_T ? _GEN_778 : _GEN_548; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_813 = _io_registerFile_2_valid_T ? _GEN_779 : _GEN_549; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_814 = _io_registerFile_2_valid_T ? _GEN_780 : _GEN_550; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_815 = _io_registerFile_2_valid_T ? _GEN_781 : _GEN_551; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_816 = _io_registerFile_2_valid_T ? _GEN_782 : _GEN_552; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_817 = _io_registerFile_2_valid_T ? _GEN_783 : _GEN_553; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_818 = _io_registerFile_2_valid_T ? _GEN_784 : _GEN_554; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_819 = _io_registerFile_2_valid_T ? _GEN_785 : _GEN_555; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_820 = _io_registerFile_2_valid_T ? _GEN_786 : _GEN_556; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_821 = _io_registerFile_2_valid_T ? _GEN_787 : _GEN_557; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_822 = _io_registerFile_2_valid_T ? _GEN_788 : _GEN_558; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_823 = _io_registerFile_2_valid_T ? _GEN_789 : _GEN_559; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_824 = _io_registerFile_2_valid_T ? _GEN_790 : _GEN_560; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_825 = _io_registerFile_2_valid_T ? _GEN_791 : _GEN_561; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_826 = _io_registerFile_2_valid_T ? _GEN_792 : _GEN_562; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_827 = _io_registerFile_2_valid_T ? _GEN_793 : _GEN_563; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_828 = _io_registerFile_2_valid_T ? _GEN_794 : _GEN_564; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_829 = _io_registerFile_2_valid_T ? _GEN_795 : _GEN_565; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_830 = _io_registerFile_2_valid_T ? _GEN_796 : _GEN_566; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_831 = _io_registerFile_2_valid_T ? _GEN_797 : _GEN_567; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_832 = _io_registerFile_2_valid_T ? _GEN_798 : _GEN_568; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_833 = _io_registerFile_2_valid_T ? _GEN_799 : _GEN_569; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_834 = _io_registerFile_2_valid_T ? _GEN_800 : _GEN_570; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_835 = _io_registerFile_2_valid_T ? _GEN_801 : _GEN_571; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_836 = _io_registerFile_2_valid_T ? _GEN_802 : _GEN_572; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_837 = _io_registerFile_2_valid_T ? _GEN_803 : _GEN_573; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_838 = _io_registerFile_2_valid_T ? _GEN_804 : _GEN_574; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_839 = _io_registerFile_2_valid_T ? _GEN_805 : _GEN_575; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_840 = _io_registerFile_2_valid_T ? _GEN_806 : _GEN_576; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_841 = _io_registerFile_2_valid_T ? _GEN_807 : _GEN_577; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_844 = _io_registerFile_2_valid_T ? _GEN_580 : 1'h1; // @[ReorderBuffer.scala 102:20 89:22]
  wire  _GEN_848 = canCommit_2 ? _GEN_811 : _GEN_547; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_849 = canCommit_2 ? _GEN_812 : _GEN_548; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_850 = canCommit_2 ? _GEN_813 : _GEN_549; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_851 = canCommit_2 ? _GEN_814 : _GEN_550; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_852 = canCommit_2 ? _GEN_815 : _GEN_551; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_853 = canCommit_2 ? _GEN_816 : _GEN_552; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_854 = canCommit_2 ? _GEN_817 : _GEN_553; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_855 = canCommit_2 ? _GEN_818 : _GEN_554; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_856 = canCommit_2 ? _GEN_819 : _GEN_555; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_857 = canCommit_2 ? _GEN_820 : _GEN_556; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_858 = canCommit_2 ? _GEN_821 : _GEN_557; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_859 = canCommit_2 ? _GEN_822 : _GEN_558; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_860 = canCommit_2 ? _GEN_823 : _GEN_559; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_861 = canCommit_2 ? _GEN_824 : _GEN_560; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_862 = canCommit_2 ? _GEN_825 : _GEN_561; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_863 = canCommit_2 ? _GEN_826 : _GEN_562; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_864 = canCommit_2 ? _GEN_827 : _GEN_563; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_865 = canCommit_2 ? _GEN_828 : _GEN_564; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_866 = canCommit_2 ? _GEN_829 : _GEN_565; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_867 = canCommit_2 ? _GEN_830 : _GEN_566; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_868 = canCommit_2 ? _GEN_831 : _GEN_567; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_869 = canCommit_2 ? _GEN_832 : _GEN_568; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_870 = canCommit_2 ? _GEN_833 : _GEN_569; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_871 = canCommit_2 ? _GEN_834 : _GEN_570; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_872 = canCommit_2 ? _GEN_835 : _GEN_571; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_873 = canCommit_2 ? _GEN_836 : _GEN_572; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_874 = canCommit_2 ? _GEN_837 : _GEN_573; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_875 = canCommit_2 ? _GEN_838 : _GEN_574; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_876 = canCommit_2 ? _GEN_839 : _GEN_575; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_877 = canCommit_2 ? _GEN_840 : _GEN_576; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_878 = canCommit_2 ? _GEN_841 : _GEN_577; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_881 = canCommit_2 ? _GEN_844 : _GEN_580; // @[ReorderBuffer.scala 88:21]
  wire [3:0] index_3 = tail + 4'h3; // @[ReorderBuffer.scala 77:22]
  wire  _GEN_902 = 4'h1 == index_3 ? buffer_1_valueReady : buffer_0_valueReady; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_903 = 4'h2 == index_3 ? buffer_2_valueReady : _GEN_902; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_904 = 4'h3 == index_3 ? buffer_3_valueReady : _GEN_903; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_905 = 4'h4 == index_3 ? buffer_4_valueReady : _GEN_904; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_906 = 4'h5 == index_3 ? buffer_5_valueReady : _GEN_905; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_907 = 4'h6 == index_3 ? buffer_6_valueReady : _GEN_906; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_908 = 4'h7 == index_3 ? buffer_7_valueReady : _GEN_907; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_909 = 4'h8 == index_3 ? buffer_8_valueReady : _GEN_908; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_910 = 4'h9 == index_3 ? buffer_9_valueReady : _GEN_909; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_911 = 4'ha == index_3 ? buffer_10_valueReady : _GEN_910; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_912 = 4'hb == index_3 ? buffer_11_valueReady : _GEN_911; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_913 = 4'hc == index_3 ? buffer_12_valueReady : _GEN_912; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_914 = 4'hd == index_3 ? buffer_13_valueReady : _GEN_913; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_915 = 4'he == index_3 ? buffer_14_valueReady : _GEN_914; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_916 = 4'hf == index_3 ? buffer_15_valueReady : _GEN_915; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_918 = 4'h1 == index_3 ? buffer_1_storeSign : buffer_0_storeSign; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_919 = 4'h2 == index_3 ? buffer_2_storeSign : _GEN_918; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_920 = 4'h3 == index_3 ? buffer_3_storeSign : _GEN_919; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_921 = 4'h4 == index_3 ? buffer_4_storeSign : _GEN_920; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_922 = 4'h5 == index_3 ? buffer_5_storeSign : _GEN_921; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_923 = 4'h6 == index_3 ? buffer_6_storeSign : _GEN_922; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_924 = 4'h7 == index_3 ? buffer_7_storeSign : _GEN_923; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_925 = 4'h8 == index_3 ? buffer_8_storeSign : _GEN_924; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_926 = 4'h9 == index_3 ? buffer_9_storeSign : _GEN_925; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_927 = 4'ha == index_3 ? buffer_10_storeSign : _GEN_926; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_928 = 4'hb == index_3 ? buffer_11_storeSign : _GEN_927; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_929 = 4'hc == index_3 ? buffer_12_storeSign : _GEN_928; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_930 = 4'hd == index_3 ? buffer_13_storeSign : _GEN_929; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_931 = 4'he == index_3 ? buffer_14_storeSign : _GEN_930; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_932 = 4'hf == index_3 ? buffer_15_storeSign : _GEN_931; // @[ReorderBuffer.scala 79:{50,50}]
  wire  instructionOk_3 = _GEN_916 | _GEN_932; // @[ReorderBuffer.scala 79:50]
  wire  canCommit_3 = canCommit_2 & index_3 != head & instructionOk_3; // @[ReorderBuffer.scala 80:49]
  wire  _GEN_934 = 4'h1 == index_3 ? buffer_1_isError : buffer_0_isError; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_935 = 4'h2 == index_3 ? buffer_2_isError : _GEN_934; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_936 = 4'h3 == index_3 ? buffer_3_isError : _GEN_935; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_937 = 4'h4 == index_3 ? buffer_4_isError : _GEN_936; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_938 = 4'h5 == index_3 ? buffer_5_isError : _GEN_937; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_939 = 4'h6 == index_3 ? buffer_6_isError : _GEN_938; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_940 = 4'h7 == index_3 ? buffer_7_isError : _GEN_939; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_941 = 4'h8 == index_3 ? buffer_8_isError : _GEN_940; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_942 = 4'h9 == index_3 ? buffer_9_isError : _GEN_941; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_943 = 4'ha == index_3 ? buffer_10_isError : _GEN_942; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_944 = 4'hb == index_3 ? buffer_11_isError : _GEN_943; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_945 = 4'hc == index_3 ? buffer_12_isError : _GEN_944; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_946 = 4'hd == index_3 ? buffer_13_isError : _GEN_945; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_947 = 4'he == index_3 ? buffer_14_isError : _GEN_946; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_948 = 4'hf == index_3 ? buffer_15_isError : _GEN_947; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _io_registerFile_3_valid_T = ~_GEN_948; // @[ReorderBuffer.scala 83:30]
  wire [63:0] _GEN_950 = 4'h1 == index_3 ? buffer_1_value : buffer_0_value; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_951 = 4'h2 == index_3 ? buffer_2_value : _GEN_950; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_952 = 4'h3 == index_3 ? buffer_3_value : _GEN_951; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_953 = 4'h4 == index_3 ? buffer_4_value : _GEN_952; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_954 = 4'h5 == index_3 ? buffer_5_value : _GEN_953; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_955 = 4'h6 == index_3 ? buffer_6_value : _GEN_954; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_956 = 4'h7 == index_3 ? buffer_7_value : _GEN_955; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_957 = 4'h8 == index_3 ? buffer_8_value : _GEN_956; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_958 = 4'h9 == index_3 ? buffer_9_value : _GEN_957; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_959 = 4'ha == index_3 ? buffer_10_value : _GEN_958; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_960 = 4'hb == index_3 ? buffer_11_value : _GEN_959; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_961 = 4'hc == index_3 ? buffer_12_value : _GEN_960; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_962 = 4'hd == index_3 ? buffer_13_value : _GEN_961; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_963 = 4'he == index_3 ? buffer_14_value : _GEN_962; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_964 = 4'hf == index_3 ? buffer_15_value : _GEN_963; // @[ReorderBuffer.scala 90:{23,23}]
  wire [4:0] _GEN_966 = 4'h1 == index_3 ? buffer_1_destinationRegister : buffer_0_destinationRegister; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_967 = 4'h2 == index_3 ? buffer_2_destinationRegister : _GEN_966; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_968 = 4'h3 == index_3 ? buffer_3_destinationRegister : _GEN_967; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_969 = 4'h4 == index_3 ? buffer_4_destinationRegister : _GEN_968; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_970 = 4'h5 == index_3 ? buffer_5_destinationRegister : _GEN_969; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_971 = 4'h6 == index_3 ? buffer_6_destinationRegister : _GEN_970; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_972 = 4'h7 == index_3 ? buffer_7_destinationRegister : _GEN_971; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_973 = 4'h8 == index_3 ? buffer_8_destinationRegister : _GEN_972; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_974 = 4'h9 == index_3 ? buffer_9_destinationRegister : _GEN_973; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_975 = 4'ha == index_3 ? buffer_10_destinationRegister : _GEN_974; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_976 = 4'hb == index_3 ? buffer_11_destinationRegister : _GEN_975; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_977 = 4'hc == index_3 ? buffer_12_destinationRegister : _GEN_976; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_978 = 4'hd == index_3 ? buffer_13_destinationRegister : _GEN_977; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_979 = 4'he == index_3 ? buffer_14_destinationRegister : _GEN_978; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_980 = 4'hf == index_3 ? buffer_15_destinationRegister : _GEN_979; // @[ReorderBuffer.scala 91:{37,37}]
  wire [3:0] _GEN_982 = 5'h1 == _GEN_980 ? registerTagMap_1_tagId : 4'h0; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_983 = 5'h2 == _GEN_980 ? registerTagMap_2_tagId : _GEN_982; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_984 = 5'h3 == _GEN_980 ? registerTagMap_3_tagId : _GEN_983; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_985 = 5'h4 == _GEN_980 ? registerTagMap_4_tagId : _GEN_984; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_986 = 5'h5 == _GEN_980 ? registerTagMap_5_tagId : _GEN_985; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_987 = 5'h6 == _GEN_980 ? registerTagMap_6_tagId : _GEN_986; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_988 = 5'h7 == _GEN_980 ? registerTagMap_7_tagId : _GEN_987; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_989 = 5'h8 == _GEN_980 ? registerTagMap_8_tagId : _GEN_988; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_990 = 5'h9 == _GEN_980 ? registerTagMap_9_tagId : _GEN_989; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_991 = 5'ha == _GEN_980 ? registerTagMap_10_tagId : _GEN_990; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_992 = 5'hb == _GEN_980 ? registerTagMap_11_tagId : _GEN_991; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_993 = 5'hc == _GEN_980 ? registerTagMap_12_tagId : _GEN_992; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_994 = 5'hd == _GEN_980 ? registerTagMap_13_tagId : _GEN_993; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_995 = 5'he == _GEN_980 ? registerTagMap_14_tagId : _GEN_994; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_996 = 5'hf == _GEN_980 ? registerTagMap_15_tagId : _GEN_995; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_997 = 5'h10 == _GEN_980 ? registerTagMap_16_tagId : _GEN_996; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_998 = 5'h11 == _GEN_980 ? registerTagMap_17_tagId : _GEN_997; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_999 = 5'h12 == _GEN_980 ? registerTagMap_18_tagId : _GEN_998; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_1000 = 5'h13 == _GEN_980 ? registerTagMap_19_tagId : _GEN_999; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_1001 = 5'h14 == _GEN_980 ? registerTagMap_20_tagId : _GEN_1000; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_1002 = 5'h15 == _GEN_980 ? registerTagMap_21_tagId : _GEN_1001; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_1003 = 5'h16 == _GEN_980 ? registerTagMap_22_tagId : _GEN_1002; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_1004 = 5'h17 == _GEN_980 ? registerTagMap_23_tagId : _GEN_1003; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_1005 = 5'h18 == _GEN_980 ? registerTagMap_24_tagId : _GEN_1004; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_1006 = 5'h19 == _GEN_980 ? registerTagMap_25_tagId : _GEN_1005; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_1007 = 5'h1a == _GEN_980 ? registerTagMap_26_tagId : _GEN_1006; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_1008 = 5'h1b == _GEN_980 ? registerTagMap_27_tagId : _GEN_1007; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_1009 = 5'h1c == _GEN_980 ? registerTagMap_28_tagId : _GEN_1008; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_1010 = 5'h1d == _GEN_980 ? registerTagMap_29_tagId : _GEN_1009; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_1011 = 5'h1e == _GEN_980 ? registerTagMap_30_tagId : _GEN_1010; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_1012 = 5'h1f == _GEN_980 ? registerTagMap_31_tagId : _GEN_1011; // @[ReorderBuffer.scala 93:{17,17}]
  wire  _T_7 = index_3 == _GEN_1012; // @[ReorderBuffer.scala 93:17]
  wire  _GEN_1046 = 5'h1 == _GEN_980 ? 1'h0 : _GEN_848; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_1047 = 5'h2 == _GEN_980 ? 1'h0 : _GEN_849; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_1048 = 5'h3 == _GEN_980 ? 1'h0 : _GEN_850; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_1049 = 5'h4 == _GEN_980 ? 1'h0 : _GEN_851; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_1050 = 5'h5 == _GEN_980 ? 1'h0 : _GEN_852; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_1051 = 5'h6 == _GEN_980 ? 1'h0 : _GEN_853; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_1052 = 5'h7 == _GEN_980 ? 1'h0 : _GEN_854; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_1053 = 5'h8 == _GEN_980 ? 1'h0 : _GEN_855; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_1054 = 5'h9 == _GEN_980 ? 1'h0 : _GEN_856; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_1055 = 5'ha == _GEN_980 ? 1'h0 : _GEN_857; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_1056 = 5'hb == _GEN_980 ? 1'h0 : _GEN_858; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_1057 = 5'hc == _GEN_980 ? 1'h0 : _GEN_859; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_1058 = 5'hd == _GEN_980 ? 1'h0 : _GEN_860; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_1059 = 5'he == _GEN_980 ? 1'h0 : _GEN_861; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_1060 = 5'hf == _GEN_980 ? 1'h0 : _GEN_862; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_1061 = 5'h10 == _GEN_980 ? 1'h0 : _GEN_863; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_1062 = 5'h11 == _GEN_980 ? 1'h0 : _GEN_864; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_1063 = 5'h12 == _GEN_980 ? 1'h0 : _GEN_865; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_1064 = 5'h13 == _GEN_980 ? 1'h0 : _GEN_866; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_1065 = 5'h14 == _GEN_980 ? 1'h0 : _GEN_867; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_1066 = 5'h15 == _GEN_980 ? 1'h0 : _GEN_868; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_1067 = 5'h16 == _GEN_980 ? 1'h0 : _GEN_869; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_1068 = 5'h17 == _GEN_980 ? 1'h0 : _GEN_870; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_1069 = 5'h18 == _GEN_980 ? 1'h0 : _GEN_871; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_1070 = 5'h19 == _GEN_980 ? 1'h0 : _GEN_872; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_1071 = 5'h1a == _GEN_980 ? 1'h0 : _GEN_873; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_1072 = 5'h1b == _GEN_980 ? 1'h0 : _GEN_874; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_1073 = 5'h1c == _GEN_980 ? 1'h0 : _GEN_875; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_1074 = 5'h1d == _GEN_980 ? 1'h0 : _GEN_876; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_1075 = 5'h1e == _GEN_980 ? 1'h0 : _GEN_877; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_1076 = 5'h1f == _GEN_980 ? 1'h0 : _GEN_878; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_1078 = _T_7 ? _GEN_1046 : _GEN_848; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_1079 = _T_7 ? _GEN_1047 : _GEN_849; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_1080 = _T_7 ? _GEN_1048 : _GEN_850; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_1081 = _T_7 ? _GEN_1049 : _GEN_851; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_1082 = _T_7 ? _GEN_1050 : _GEN_852; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_1083 = _T_7 ? _GEN_1051 : _GEN_853; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_1084 = _T_7 ? _GEN_1052 : _GEN_854; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_1085 = _T_7 ? _GEN_1053 : _GEN_855; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_1086 = _T_7 ? _GEN_1054 : _GEN_856; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_1087 = _T_7 ? _GEN_1055 : _GEN_857; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_1088 = _T_7 ? _GEN_1056 : _GEN_858; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_1089 = _T_7 ? _GEN_1057 : _GEN_859; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_1090 = _T_7 ? _GEN_1058 : _GEN_860; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_1091 = _T_7 ? _GEN_1059 : _GEN_861; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_1092 = _T_7 ? _GEN_1060 : _GEN_862; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_1093 = _T_7 ? _GEN_1061 : _GEN_863; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_1094 = _T_7 ? _GEN_1062 : _GEN_864; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_1095 = _T_7 ? _GEN_1063 : _GEN_865; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_1096 = _T_7 ? _GEN_1064 : _GEN_866; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_1097 = _T_7 ? _GEN_1065 : _GEN_867; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_1098 = _T_7 ? _GEN_1066 : _GEN_868; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_1099 = _T_7 ? _GEN_1067 : _GEN_869; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_1100 = _T_7 ? _GEN_1068 : _GEN_870; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_1101 = _T_7 ? _GEN_1069 : _GEN_871; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_1102 = _T_7 ? _GEN_1070 : _GEN_872; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_1103 = _T_7 ? _GEN_1071 : _GEN_873; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_1104 = _T_7 ? _GEN_1072 : _GEN_874; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_1105 = _T_7 ? _GEN_1073 : _GEN_875; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_1106 = _T_7 ? _GEN_1074 : _GEN_876; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_1107 = _T_7 ? _GEN_1075 : _GEN_877; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_1108 = _T_7 ? _GEN_1076 : _GEN_878; // @[ReorderBuffer.scala 94:11]
  wire [63:0] _GEN_1109 = _io_registerFile_3_valid_T ? _GEN_964 : 64'h0; // @[ReorderBuffer.scala 84:19 89:22 90:23]
  wire [4:0] _GEN_1110 = _io_registerFile_3_valid_T ? _GEN_980 : 5'h0; // @[ReorderBuffer.scala 89:22 85:33 91:37]
  wire  _GEN_1112 = _io_registerFile_3_valid_T ? _GEN_1078 : _GEN_848; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_1113 = _io_registerFile_3_valid_T ? _GEN_1079 : _GEN_849; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_1114 = _io_registerFile_3_valid_T ? _GEN_1080 : _GEN_850; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_1115 = _io_registerFile_3_valid_T ? _GEN_1081 : _GEN_851; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_1116 = _io_registerFile_3_valid_T ? _GEN_1082 : _GEN_852; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_1117 = _io_registerFile_3_valid_T ? _GEN_1083 : _GEN_853; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_1118 = _io_registerFile_3_valid_T ? _GEN_1084 : _GEN_854; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_1119 = _io_registerFile_3_valid_T ? _GEN_1085 : _GEN_855; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_1120 = _io_registerFile_3_valid_T ? _GEN_1086 : _GEN_856; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_1121 = _io_registerFile_3_valid_T ? _GEN_1087 : _GEN_857; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_1122 = _io_registerFile_3_valid_T ? _GEN_1088 : _GEN_858; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_1123 = _io_registerFile_3_valid_T ? _GEN_1089 : _GEN_859; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_1124 = _io_registerFile_3_valid_T ? _GEN_1090 : _GEN_860; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_1125 = _io_registerFile_3_valid_T ? _GEN_1091 : _GEN_861; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_1126 = _io_registerFile_3_valid_T ? _GEN_1092 : _GEN_862; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_1127 = _io_registerFile_3_valid_T ? _GEN_1093 : _GEN_863; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_1128 = _io_registerFile_3_valid_T ? _GEN_1094 : _GEN_864; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_1129 = _io_registerFile_3_valid_T ? _GEN_1095 : _GEN_865; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_1130 = _io_registerFile_3_valid_T ? _GEN_1096 : _GEN_866; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_1131 = _io_registerFile_3_valid_T ? _GEN_1097 : _GEN_867; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_1132 = _io_registerFile_3_valid_T ? _GEN_1098 : _GEN_868; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_1133 = _io_registerFile_3_valid_T ? _GEN_1099 : _GEN_869; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_1134 = _io_registerFile_3_valid_T ? _GEN_1100 : _GEN_870; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_1135 = _io_registerFile_3_valid_T ? _GEN_1101 : _GEN_871; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_1136 = _io_registerFile_3_valid_T ? _GEN_1102 : _GEN_872; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_1137 = _io_registerFile_3_valid_T ? _GEN_1103 : _GEN_873; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_1138 = _io_registerFile_3_valid_T ? _GEN_1104 : _GEN_874; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_1139 = _io_registerFile_3_valid_T ? _GEN_1105 : _GEN_875; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_1140 = _io_registerFile_3_valid_T ? _GEN_1106 : _GEN_876; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_1141 = _io_registerFile_3_valid_T ? _GEN_1107 : _GEN_877; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_1142 = _io_registerFile_3_valid_T ? _GEN_1108 : _GEN_878; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_1145 = _io_registerFile_3_valid_T ? _GEN_881 : 1'h1; // @[ReorderBuffer.scala 102:20 89:22]
  wire  _GEN_1149 = canCommit_3 ? _GEN_1112 : _GEN_848; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_1150 = canCommit_3 ? _GEN_1113 : _GEN_849; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_1151 = canCommit_3 ? _GEN_1114 : _GEN_850; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_1152 = canCommit_3 ? _GEN_1115 : _GEN_851; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_1153 = canCommit_3 ? _GEN_1116 : _GEN_852; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_1154 = canCommit_3 ? _GEN_1117 : _GEN_853; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_1155 = canCommit_3 ? _GEN_1118 : _GEN_854; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_1156 = canCommit_3 ? _GEN_1119 : _GEN_855; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_1157 = canCommit_3 ? _GEN_1120 : _GEN_856; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_1158 = canCommit_3 ? _GEN_1121 : _GEN_857; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_1159 = canCommit_3 ? _GEN_1122 : _GEN_858; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_1160 = canCommit_3 ? _GEN_1123 : _GEN_859; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_1161 = canCommit_3 ? _GEN_1124 : _GEN_860; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_1162 = canCommit_3 ? _GEN_1125 : _GEN_861; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_1163 = canCommit_3 ? _GEN_1126 : _GEN_862; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_1164 = canCommit_3 ? _GEN_1127 : _GEN_863; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_1165 = canCommit_3 ? _GEN_1128 : _GEN_864; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_1166 = canCommit_3 ? _GEN_1129 : _GEN_865; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_1167 = canCommit_3 ? _GEN_1130 : _GEN_866; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_1168 = canCommit_3 ? _GEN_1131 : _GEN_867; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_1169 = canCommit_3 ? _GEN_1132 : _GEN_868; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_1170 = canCommit_3 ? _GEN_1133 : _GEN_869; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_1171 = canCommit_3 ? _GEN_1134 : _GEN_870; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_1172 = canCommit_3 ? _GEN_1135 : _GEN_871; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_1173 = canCommit_3 ? _GEN_1136 : _GEN_872; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_1174 = canCommit_3 ? _GEN_1137 : _GEN_873; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_1175 = canCommit_3 ? _GEN_1138 : _GEN_874; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_1176 = canCommit_3 ? _GEN_1139 : _GEN_875; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_1177 = canCommit_3 ? _GEN_1140 : _GEN_876; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_1178 = canCommit_3 ? _GEN_1141 : _GEN_877; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_1179 = canCommit_3 ? _GEN_1142 : _GEN_878; // @[ReorderBuffer.scala 88:21]
  wire  _tailDelta_T = ~io_registerFile_0_valid; // @[ReorderBuffer.scala 120:7]
  wire  _tailDelta_T_1 = ~io_registerFile_1_valid; // @[ReorderBuffer.scala 120:7]
  wire  _tailDelta_T_2 = ~io_registerFile_2_valid; // @[ReorderBuffer.scala 120:7]
  wire  _tailDelta_T_3 = ~io_registerFile_3_valid; // @[ReorderBuffer.scala 120:7]
  wire [2:0] _tailDelta_T_4 = _tailDelta_T_3 ? 3'h3 : 3'h4; // @[Mux.scala 101:16]
  wire [2:0] _tailDelta_T_5 = _tailDelta_T_2 ? 3'h2 : _tailDelta_T_4; // @[Mux.scala 101:16]
  wire [2:0] _tailDelta_T_6 = _tailDelta_T_1 ? 3'h1 : _tailDelta_T_5; // @[Mux.scala 101:16]
  wire [2:0] tailDelta = _tailDelta_T ? 3'h0 : _tailDelta_T_6; // @[Mux.scala 101:16]
  wire [3:0] _io_decoders_0_ready_T_1 = head + 4'h1; // @[ReorderBuffer.scala 129:48]
  wire  _T_8 = io_decoders_0_valid & io_decoders_0_ready; // @[ReorderBuffer.scala 130:24]
  wire  _GEN_1218 = 4'h0 == head ? 1'h0 : buffer_0_valueReady; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire  _GEN_1219 = 4'h1 == head ? 1'h0 : buffer_1_valueReady; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire  _GEN_1220 = 4'h2 == head ? 1'h0 : buffer_2_valueReady; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire  _GEN_1221 = 4'h3 == head ? 1'h0 : buffer_3_valueReady; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire  _GEN_1222 = 4'h4 == head ? 1'h0 : buffer_4_valueReady; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire  _GEN_1223 = 4'h5 == head ? 1'h0 : buffer_5_valueReady; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire  _GEN_1224 = 4'h6 == head ? 1'h0 : buffer_6_valueReady; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire  _GEN_1225 = 4'h7 == head ? 1'h0 : buffer_7_valueReady; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire  _GEN_1226 = 4'h8 == head ? 1'h0 : buffer_8_valueReady; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire  _GEN_1227 = 4'h9 == head ? 1'h0 : buffer_9_valueReady; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire  _GEN_1228 = 4'ha == head ? 1'h0 : buffer_10_valueReady; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire  _GEN_1229 = 4'hb == head ? 1'h0 : buffer_11_valueReady; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire  _GEN_1230 = 4'hc == head ? 1'h0 : buffer_12_valueReady; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire  _GEN_1231 = 4'hd == head ? 1'h0 : buffer_13_valueReady; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire  _GEN_1232 = 4'he == head ? 1'h0 : buffer_14_valueReady; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire  _GEN_1233 = 4'hf == head ? 1'h0 : buffer_15_valueReady; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire [63:0] _GEN_1234 = 4'h0 == head ? 64'h0 : buffer_0_value; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire [63:0] _GEN_1235 = 4'h1 == head ? 64'h0 : buffer_1_value; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire [63:0] _GEN_1236 = 4'h2 == head ? 64'h0 : buffer_2_value; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire [63:0] _GEN_1237 = 4'h3 == head ? 64'h0 : buffer_3_value; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire [63:0] _GEN_1238 = 4'h4 == head ? 64'h0 : buffer_4_value; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire [63:0] _GEN_1239 = 4'h5 == head ? 64'h0 : buffer_5_value; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire [63:0] _GEN_1240 = 4'h6 == head ? 64'h0 : buffer_6_value; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire [63:0] _GEN_1241 = 4'h7 == head ? 64'h0 : buffer_7_value; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire [63:0] _GEN_1242 = 4'h8 == head ? 64'h0 : buffer_8_value; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire [63:0] _GEN_1243 = 4'h9 == head ? 64'h0 : buffer_9_value; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire [63:0] _GEN_1244 = 4'ha == head ? 64'h0 : buffer_10_value; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire [63:0] _GEN_1245 = 4'hb == head ? 64'h0 : buffer_11_value; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire [63:0] _GEN_1246 = 4'hc == head ? 64'h0 : buffer_12_value; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire [63:0] _GEN_1247 = 4'hd == head ? 64'h0 : buffer_13_value; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire [63:0] _GEN_1248 = 4'he == head ? 64'h0 : buffer_14_value; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire [63:0] _GEN_1249 = 4'hf == head ? 64'h0 : buffer_15_value; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire  _GEN_1282 = 4'h0 == head ? 1'h0 : buffer_0_isError; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire  _GEN_1283 = 4'h1 == head ? 1'h0 : buffer_1_isError; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire  _GEN_1284 = 4'h2 == head ? 1'h0 : buffer_2_isError; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire  _GEN_1285 = 4'h3 == head ? 1'h0 : buffer_3_isError; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire  _GEN_1286 = 4'h4 == head ? 1'h0 : buffer_4_isError; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire  _GEN_1287 = 4'h5 == head ? 1'h0 : buffer_5_isError; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire  _GEN_1288 = 4'h6 == head ? 1'h0 : buffer_6_isError; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire  _GEN_1289 = 4'h7 == head ? 1'h0 : buffer_7_isError; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire  _GEN_1290 = 4'h8 == head ? 1'h0 : buffer_8_isError; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire  _GEN_1291 = 4'h9 == head ? 1'h0 : buffer_9_isError; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire  _GEN_1292 = 4'ha == head ? 1'h0 : buffer_10_isError; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire  _GEN_1293 = 4'hb == head ? 1'h0 : buffer_11_isError; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire  _GEN_1294 = 4'hc == head ? 1'h0 : buffer_12_isError; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire  _GEN_1295 = 4'hd == head ? 1'h0 : buffer_13_isError; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire  _GEN_1296 = 4'he == head ? 1'h0 : buffer_14_isError; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire  _GEN_1297 = 4'hf == head ? 1'h0 : buffer_15_isError; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire  _GEN_1314 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1218 : buffer_0_valueReady; // @[ReorderBuffer.scala 130:42 55:23]
  wire  _GEN_1315 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1219 : buffer_1_valueReady; // @[ReorderBuffer.scala 130:42 55:23]
  wire  _GEN_1316 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1220 : buffer_2_valueReady; // @[ReorderBuffer.scala 130:42 55:23]
  wire  _GEN_1317 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1221 : buffer_3_valueReady; // @[ReorderBuffer.scala 130:42 55:23]
  wire  _GEN_1318 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1222 : buffer_4_valueReady; // @[ReorderBuffer.scala 130:42 55:23]
  wire  _GEN_1319 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1223 : buffer_5_valueReady; // @[ReorderBuffer.scala 130:42 55:23]
  wire  _GEN_1320 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1224 : buffer_6_valueReady; // @[ReorderBuffer.scala 130:42 55:23]
  wire  _GEN_1321 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1225 : buffer_7_valueReady; // @[ReorderBuffer.scala 130:42 55:23]
  wire  _GEN_1322 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1226 : buffer_8_valueReady; // @[ReorderBuffer.scala 130:42 55:23]
  wire  _GEN_1323 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1227 : buffer_9_valueReady; // @[ReorderBuffer.scala 130:42 55:23]
  wire  _GEN_1324 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1228 : buffer_10_valueReady; // @[ReorderBuffer.scala 130:42 55:23]
  wire  _GEN_1325 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1229 : buffer_11_valueReady; // @[ReorderBuffer.scala 130:42 55:23]
  wire  _GEN_1326 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1230 : buffer_12_valueReady; // @[ReorderBuffer.scala 130:42 55:23]
  wire  _GEN_1327 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1231 : buffer_13_valueReady; // @[ReorderBuffer.scala 130:42 55:23]
  wire  _GEN_1328 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1232 : buffer_14_valueReady; // @[ReorderBuffer.scala 130:42 55:23]
  wire  _GEN_1329 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1233 : buffer_15_valueReady; // @[ReorderBuffer.scala 130:42 55:23]
  wire [63:0] _GEN_1330 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1234 : buffer_0_value; // @[ReorderBuffer.scala 130:42 55:23]
  wire [63:0] _GEN_1331 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1235 : buffer_1_value; // @[ReorderBuffer.scala 130:42 55:23]
  wire [63:0] _GEN_1332 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1236 : buffer_2_value; // @[ReorderBuffer.scala 130:42 55:23]
  wire [63:0] _GEN_1333 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1237 : buffer_3_value; // @[ReorderBuffer.scala 130:42 55:23]
  wire [63:0] _GEN_1334 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1238 : buffer_4_value; // @[ReorderBuffer.scala 130:42 55:23]
  wire [63:0] _GEN_1335 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1239 : buffer_5_value; // @[ReorderBuffer.scala 130:42 55:23]
  wire [63:0] _GEN_1336 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1240 : buffer_6_value; // @[ReorderBuffer.scala 130:42 55:23]
  wire [63:0] _GEN_1337 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1241 : buffer_7_value; // @[ReorderBuffer.scala 130:42 55:23]
  wire [63:0] _GEN_1338 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1242 : buffer_8_value; // @[ReorderBuffer.scala 130:42 55:23]
  wire [63:0] _GEN_1339 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1243 : buffer_9_value; // @[ReorderBuffer.scala 130:42 55:23]
  wire [63:0] _GEN_1340 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1244 : buffer_10_value; // @[ReorderBuffer.scala 130:42 55:23]
  wire [63:0] _GEN_1341 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1245 : buffer_11_value; // @[ReorderBuffer.scala 130:42 55:23]
  wire [63:0] _GEN_1342 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1246 : buffer_12_value; // @[ReorderBuffer.scala 130:42 55:23]
  wire [63:0] _GEN_1343 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1247 : buffer_13_value; // @[ReorderBuffer.scala 130:42 55:23]
  wire [63:0] _GEN_1344 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1248 : buffer_14_value; // @[ReorderBuffer.scala 130:42 55:23]
  wire [63:0] _GEN_1345 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1249 : buffer_15_value; // @[ReorderBuffer.scala 130:42 55:23]
  wire  _GEN_1378 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1282 : buffer_0_isError; // @[ReorderBuffer.scala 130:42 55:23]
  wire  _GEN_1379 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1283 : buffer_1_isError; // @[ReorderBuffer.scala 130:42 55:23]
  wire  _GEN_1380 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1284 : buffer_2_isError; // @[ReorderBuffer.scala 130:42 55:23]
  wire  _GEN_1381 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1285 : buffer_3_isError; // @[ReorderBuffer.scala 130:42 55:23]
  wire  _GEN_1382 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1286 : buffer_4_isError; // @[ReorderBuffer.scala 130:42 55:23]
  wire  _GEN_1383 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1287 : buffer_5_isError; // @[ReorderBuffer.scala 130:42 55:23]
  wire  _GEN_1384 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1288 : buffer_6_isError; // @[ReorderBuffer.scala 130:42 55:23]
  wire  _GEN_1385 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1289 : buffer_7_isError; // @[ReorderBuffer.scala 130:42 55:23]
  wire  _GEN_1386 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1290 : buffer_8_isError; // @[ReorderBuffer.scala 130:42 55:23]
  wire  _GEN_1387 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1291 : buffer_9_isError; // @[ReorderBuffer.scala 130:42 55:23]
  wire  _GEN_1388 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1292 : buffer_10_isError; // @[ReorderBuffer.scala 130:42 55:23]
  wire  _GEN_1389 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1293 : buffer_11_isError; // @[ReorderBuffer.scala 130:42 55:23]
  wire  _GEN_1390 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1294 : buffer_12_isError; // @[ReorderBuffer.scala 130:42 55:23]
  wire  _GEN_1391 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1295 : buffer_13_isError; // @[ReorderBuffer.scala 130:42 55:23]
  wire  _GEN_1392 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1296 : buffer_14_isError; // @[ReorderBuffer.scala 130:42 55:23]
  wire  _GEN_1393 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1297 : buffer_15_isError; // @[ReorderBuffer.scala 130:42 55:23]
  wire  _GEN_1395 = 5'h1 == io_decoders_0_destination_destinationRegister | _GEN_1149; // @[ReorderBuffer.scala 146:{69,69}]
  wire  _GEN_1396 = 5'h2 == io_decoders_0_destination_destinationRegister | _GEN_1150; // @[ReorderBuffer.scala 146:{69,69}]
  wire  _GEN_1397 = 5'h3 == io_decoders_0_destination_destinationRegister | _GEN_1151; // @[ReorderBuffer.scala 146:{69,69}]
  wire  _GEN_1398 = 5'h4 == io_decoders_0_destination_destinationRegister | _GEN_1152; // @[ReorderBuffer.scala 146:{69,69}]
  wire  _GEN_1399 = 5'h5 == io_decoders_0_destination_destinationRegister | _GEN_1153; // @[ReorderBuffer.scala 146:{69,69}]
  wire  _GEN_1400 = 5'h6 == io_decoders_0_destination_destinationRegister | _GEN_1154; // @[ReorderBuffer.scala 146:{69,69}]
  wire  _GEN_1401 = 5'h7 == io_decoders_0_destination_destinationRegister | _GEN_1155; // @[ReorderBuffer.scala 146:{69,69}]
  wire  _GEN_1402 = 5'h8 == io_decoders_0_destination_destinationRegister | _GEN_1156; // @[ReorderBuffer.scala 146:{69,69}]
  wire  _GEN_1403 = 5'h9 == io_decoders_0_destination_destinationRegister | _GEN_1157; // @[ReorderBuffer.scala 146:{69,69}]
  wire  _GEN_1404 = 5'ha == io_decoders_0_destination_destinationRegister | _GEN_1158; // @[ReorderBuffer.scala 146:{69,69}]
  wire  _GEN_1405 = 5'hb == io_decoders_0_destination_destinationRegister | _GEN_1159; // @[ReorderBuffer.scala 146:{69,69}]
  wire  _GEN_1406 = 5'hc == io_decoders_0_destination_destinationRegister | _GEN_1160; // @[ReorderBuffer.scala 146:{69,69}]
  wire  _GEN_1407 = 5'hd == io_decoders_0_destination_destinationRegister | _GEN_1161; // @[ReorderBuffer.scala 146:{69,69}]
  wire  _GEN_1408 = 5'he == io_decoders_0_destination_destinationRegister | _GEN_1162; // @[ReorderBuffer.scala 146:{69,69}]
  wire  _GEN_1409 = 5'hf == io_decoders_0_destination_destinationRegister | _GEN_1163; // @[ReorderBuffer.scala 146:{69,69}]
  wire  _GEN_1410 = 5'h10 == io_decoders_0_destination_destinationRegister | _GEN_1164; // @[ReorderBuffer.scala 146:{69,69}]
  wire  _GEN_1411 = 5'h11 == io_decoders_0_destination_destinationRegister | _GEN_1165; // @[ReorderBuffer.scala 146:{69,69}]
  wire  _GEN_1412 = 5'h12 == io_decoders_0_destination_destinationRegister | _GEN_1166; // @[ReorderBuffer.scala 146:{69,69}]
  wire  _GEN_1413 = 5'h13 == io_decoders_0_destination_destinationRegister | _GEN_1167; // @[ReorderBuffer.scala 146:{69,69}]
  wire  _GEN_1414 = 5'h14 == io_decoders_0_destination_destinationRegister | _GEN_1168; // @[ReorderBuffer.scala 146:{69,69}]
  wire  _GEN_1415 = 5'h15 == io_decoders_0_destination_destinationRegister | _GEN_1169; // @[ReorderBuffer.scala 146:{69,69}]
  wire  _GEN_1416 = 5'h16 == io_decoders_0_destination_destinationRegister | _GEN_1170; // @[ReorderBuffer.scala 146:{69,69}]
  wire  _GEN_1417 = 5'h17 == io_decoders_0_destination_destinationRegister | _GEN_1171; // @[ReorderBuffer.scala 146:{69,69}]
  wire  _GEN_1418 = 5'h18 == io_decoders_0_destination_destinationRegister | _GEN_1172; // @[ReorderBuffer.scala 146:{69,69}]
  wire  _GEN_1419 = 5'h19 == io_decoders_0_destination_destinationRegister | _GEN_1173; // @[ReorderBuffer.scala 146:{69,69}]
  wire  _GEN_1420 = 5'h1a == io_decoders_0_destination_destinationRegister | _GEN_1174; // @[ReorderBuffer.scala 146:{69,69}]
  wire  _GEN_1421 = 5'h1b == io_decoders_0_destination_destinationRegister | _GEN_1175; // @[ReorderBuffer.scala 146:{69,69}]
  wire  _GEN_1422 = 5'h1c == io_decoders_0_destination_destinationRegister | _GEN_1176; // @[ReorderBuffer.scala 146:{69,69}]
  wire  _GEN_1423 = 5'h1d == io_decoders_0_destination_destinationRegister | _GEN_1177; // @[ReorderBuffer.scala 146:{69,69}]
  wire  _GEN_1424 = 5'h1e == io_decoders_0_destination_destinationRegister | _GEN_1178; // @[ReorderBuffer.scala 146:{69,69}]
  wire  _GEN_1425 = 5'h1f == io_decoders_0_destination_destinationRegister | _GEN_1179; // @[ReorderBuffer.scala 146:{69,69}]
  wire  _GEN_1524 = 5'h2 == io_decoders_0_source1_sourceRegister ? registerTagMap_2_valid : 5'h1 ==
    io_decoders_0_source1_sourceRegister & registerTagMap_1_valid; // @[ReorderBuffer.scala 155:{41,41}]
  wire  _GEN_1525 = 5'h3 == io_decoders_0_source1_sourceRegister ? registerTagMap_3_valid : _GEN_1524; // @[ReorderBuffer.scala 155:{41,41}]
  wire  _GEN_1526 = 5'h4 == io_decoders_0_source1_sourceRegister ? registerTagMap_4_valid : _GEN_1525; // @[ReorderBuffer.scala 155:{41,41}]
  wire  _GEN_1527 = 5'h5 == io_decoders_0_source1_sourceRegister ? registerTagMap_5_valid : _GEN_1526; // @[ReorderBuffer.scala 155:{41,41}]
  wire  _GEN_1528 = 5'h6 == io_decoders_0_source1_sourceRegister ? registerTagMap_6_valid : _GEN_1527; // @[ReorderBuffer.scala 155:{41,41}]
  wire  _GEN_1529 = 5'h7 == io_decoders_0_source1_sourceRegister ? registerTagMap_7_valid : _GEN_1528; // @[ReorderBuffer.scala 155:{41,41}]
  wire  _GEN_1530 = 5'h8 == io_decoders_0_source1_sourceRegister ? registerTagMap_8_valid : _GEN_1529; // @[ReorderBuffer.scala 155:{41,41}]
  wire  _GEN_1531 = 5'h9 == io_decoders_0_source1_sourceRegister ? registerTagMap_9_valid : _GEN_1530; // @[ReorderBuffer.scala 155:{41,41}]
  wire  _GEN_1532 = 5'ha == io_decoders_0_source1_sourceRegister ? registerTagMap_10_valid : _GEN_1531; // @[ReorderBuffer.scala 155:{41,41}]
  wire  _GEN_1533 = 5'hb == io_decoders_0_source1_sourceRegister ? registerTagMap_11_valid : _GEN_1532; // @[ReorderBuffer.scala 155:{41,41}]
  wire  _GEN_1534 = 5'hc == io_decoders_0_source1_sourceRegister ? registerTagMap_12_valid : _GEN_1533; // @[ReorderBuffer.scala 155:{41,41}]
  wire  _GEN_1535 = 5'hd == io_decoders_0_source1_sourceRegister ? registerTagMap_13_valid : _GEN_1534; // @[ReorderBuffer.scala 155:{41,41}]
  wire  _GEN_1536 = 5'he == io_decoders_0_source1_sourceRegister ? registerTagMap_14_valid : _GEN_1535; // @[ReorderBuffer.scala 155:{41,41}]
  wire  _GEN_1537 = 5'hf == io_decoders_0_source1_sourceRegister ? registerTagMap_15_valid : _GEN_1536; // @[ReorderBuffer.scala 155:{41,41}]
  wire  _GEN_1538 = 5'h10 == io_decoders_0_source1_sourceRegister ? registerTagMap_16_valid : _GEN_1537; // @[ReorderBuffer.scala 155:{41,41}]
  wire  _GEN_1539 = 5'h11 == io_decoders_0_source1_sourceRegister ? registerTagMap_17_valid : _GEN_1538; // @[ReorderBuffer.scala 155:{41,41}]
  wire  _GEN_1540 = 5'h12 == io_decoders_0_source1_sourceRegister ? registerTagMap_18_valid : _GEN_1539; // @[ReorderBuffer.scala 155:{41,41}]
  wire  _GEN_1541 = 5'h13 == io_decoders_0_source1_sourceRegister ? registerTagMap_19_valid : _GEN_1540; // @[ReorderBuffer.scala 155:{41,41}]
  wire  _GEN_1542 = 5'h14 == io_decoders_0_source1_sourceRegister ? registerTagMap_20_valid : _GEN_1541; // @[ReorderBuffer.scala 155:{41,41}]
  wire  _GEN_1543 = 5'h15 == io_decoders_0_source1_sourceRegister ? registerTagMap_21_valid : _GEN_1542; // @[ReorderBuffer.scala 155:{41,41}]
  wire  _GEN_1544 = 5'h16 == io_decoders_0_source1_sourceRegister ? registerTagMap_22_valid : _GEN_1543; // @[ReorderBuffer.scala 155:{41,41}]
  wire  _GEN_1545 = 5'h17 == io_decoders_0_source1_sourceRegister ? registerTagMap_23_valid : _GEN_1544; // @[ReorderBuffer.scala 155:{41,41}]
  wire  _GEN_1546 = 5'h18 == io_decoders_0_source1_sourceRegister ? registerTagMap_24_valid : _GEN_1545; // @[ReorderBuffer.scala 155:{41,41}]
  wire  _GEN_1547 = 5'h19 == io_decoders_0_source1_sourceRegister ? registerTagMap_25_valid : _GEN_1546; // @[ReorderBuffer.scala 155:{41,41}]
  wire  _GEN_1548 = 5'h1a == io_decoders_0_source1_sourceRegister ? registerTagMap_26_valid : _GEN_1547; // @[ReorderBuffer.scala 155:{41,41}]
  wire  _GEN_1549 = 5'h1b == io_decoders_0_source1_sourceRegister ? registerTagMap_27_valid : _GEN_1548; // @[ReorderBuffer.scala 155:{41,41}]
  wire  _GEN_1550 = 5'h1c == io_decoders_0_source1_sourceRegister ? registerTagMap_28_valid : _GEN_1549; // @[ReorderBuffer.scala 155:{41,41}]
  wire  _GEN_1551 = 5'h1d == io_decoders_0_source1_sourceRegister ? registerTagMap_29_valid : _GEN_1550; // @[ReorderBuffer.scala 155:{41,41}]
  wire  _GEN_1552 = 5'h1e == io_decoders_0_source1_sourceRegister ? registerTagMap_30_valid : _GEN_1551; // @[ReorderBuffer.scala 155:{41,41}]
  wire  _GEN_1553 = 5'h1f == io_decoders_0_source1_sourceRegister ? registerTagMap_31_valid : _GEN_1552; // @[ReorderBuffer.scala 155:{41,41}]
  wire [3:0] _GEN_1555 = 5'h1 == io_decoders_0_source1_sourceRegister ? registerTagMap_1_tagId : 4'h0; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1556 = 5'h2 == io_decoders_0_source1_sourceRegister ? registerTagMap_2_tagId : _GEN_1555; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1557 = 5'h3 == io_decoders_0_source1_sourceRegister ? registerTagMap_3_tagId : _GEN_1556; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1558 = 5'h4 == io_decoders_0_source1_sourceRegister ? registerTagMap_4_tagId : _GEN_1557; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1559 = 5'h5 == io_decoders_0_source1_sourceRegister ? registerTagMap_5_tagId : _GEN_1558; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1560 = 5'h6 == io_decoders_0_source1_sourceRegister ? registerTagMap_6_tagId : _GEN_1559; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1561 = 5'h7 == io_decoders_0_source1_sourceRegister ? registerTagMap_7_tagId : _GEN_1560; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1562 = 5'h8 == io_decoders_0_source1_sourceRegister ? registerTagMap_8_tagId : _GEN_1561; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1563 = 5'h9 == io_decoders_0_source1_sourceRegister ? registerTagMap_9_tagId : _GEN_1562; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1564 = 5'ha == io_decoders_0_source1_sourceRegister ? registerTagMap_10_tagId : _GEN_1563; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1565 = 5'hb == io_decoders_0_source1_sourceRegister ? registerTagMap_11_tagId : _GEN_1564; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1566 = 5'hc == io_decoders_0_source1_sourceRegister ? registerTagMap_12_tagId : _GEN_1565; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1567 = 5'hd == io_decoders_0_source1_sourceRegister ? registerTagMap_13_tagId : _GEN_1566; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1568 = 5'he == io_decoders_0_source1_sourceRegister ? registerTagMap_14_tagId : _GEN_1567; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1569 = 5'hf == io_decoders_0_source1_sourceRegister ? registerTagMap_15_tagId : _GEN_1568; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1570 = 5'h10 == io_decoders_0_source1_sourceRegister ? registerTagMap_16_tagId : _GEN_1569; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1571 = 5'h11 == io_decoders_0_source1_sourceRegister ? registerTagMap_17_tagId : _GEN_1570; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1572 = 5'h12 == io_decoders_0_source1_sourceRegister ? registerTagMap_18_tagId : _GEN_1571; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1573 = 5'h13 == io_decoders_0_source1_sourceRegister ? registerTagMap_19_tagId : _GEN_1572; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1574 = 5'h14 == io_decoders_0_source1_sourceRegister ? registerTagMap_20_tagId : _GEN_1573; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1575 = 5'h15 == io_decoders_0_source1_sourceRegister ? registerTagMap_21_tagId : _GEN_1574; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1576 = 5'h16 == io_decoders_0_source1_sourceRegister ? registerTagMap_22_tagId : _GEN_1575; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1577 = 5'h17 == io_decoders_0_source1_sourceRegister ? registerTagMap_23_tagId : _GEN_1576; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1578 = 5'h18 == io_decoders_0_source1_sourceRegister ? registerTagMap_24_tagId : _GEN_1577; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1579 = 5'h19 == io_decoders_0_source1_sourceRegister ? registerTagMap_25_tagId : _GEN_1578; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1580 = 5'h1a == io_decoders_0_source1_sourceRegister ? registerTagMap_26_tagId : _GEN_1579; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1581 = 5'h1b == io_decoders_0_source1_sourceRegister ? registerTagMap_27_tagId : _GEN_1580; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1582 = 5'h1c == io_decoders_0_source1_sourceRegister ? registerTagMap_28_tagId : _GEN_1581; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1583 = 5'h1d == io_decoders_0_source1_sourceRegister ? registerTagMap_29_tagId : _GEN_1582; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1584 = 5'h1e == io_decoders_0_source1_sourceRegister ? registerTagMap_30_tagId : _GEN_1583; // @[Tag.scala 23:{10,10}]
  wire [3:0] io_decoders_0_source1_matchingTag_bits_w_id = 5'h1f == io_decoders_0_source1_sourceRegister ?
    registerTagMap_31_tagId : _GEN_1584; // @[Tag.scala 23:{10,10}]
  wire  _GEN_1587 = 4'h1 == io_decoders_0_source1_matchingTag_bits_w_id ? buffer_1_valueReady : buffer_0_valueReady; // @[ReorderBuffer.scala 160:{35,35}]
  wire  _GEN_1588 = 4'h2 == io_decoders_0_source1_matchingTag_bits_w_id ? buffer_2_valueReady : _GEN_1587; // @[ReorderBuffer.scala 160:{35,35}]
  wire  _GEN_1589 = 4'h3 == io_decoders_0_source1_matchingTag_bits_w_id ? buffer_3_valueReady : _GEN_1588; // @[ReorderBuffer.scala 160:{35,35}]
  wire  _GEN_1590 = 4'h4 == io_decoders_0_source1_matchingTag_bits_w_id ? buffer_4_valueReady : _GEN_1589; // @[ReorderBuffer.scala 160:{35,35}]
  wire  _GEN_1591 = 4'h5 == io_decoders_0_source1_matchingTag_bits_w_id ? buffer_5_valueReady : _GEN_1590; // @[ReorderBuffer.scala 160:{35,35}]
  wire  _GEN_1592 = 4'h6 == io_decoders_0_source1_matchingTag_bits_w_id ? buffer_6_valueReady : _GEN_1591; // @[ReorderBuffer.scala 160:{35,35}]
  wire  _GEN_1593 = 4'h7 == io_decoders_0_source1_matchingTag_bits_w_id ? buffer_7_valueReady : _GEN_1592; // @[ReorderBuffer.scala 160:{35,35}]
  wire  _GEN_1594 = 4'h8 == io_decoders_0_source1_matchingTag_bits_w_id ? buffer_8_valueReady : _GEN_1593; // @[ReorderBuffer.scala 160:{35,35}]
  wire  _GEN_1595 = 4'h9 == io_decoders_0_source1_matchingTag_bits_w_id ? buffer_9_valueReady : _GEN_1594; // @[ReorderBuffer.scala 160:{35,35}]
  wire  _GEN_1596 = 4'ha == io_decoders_0_source1_matchingTag_bits_w_id ? buffer_10_valueReady : _GEN_1595; // @[ReorderBuffer.scala 160:{35,35}]
  wire  _GEN_1597 = 4'hb == io_decoders_0_source1_matchingTag_bits_w_id ? buffer_11_valueReady : _GEN_1596; // @[ReorderBuffer.scala 160:{35,35}]
  wire  _GEN_1598 = 4'hc == io_decoders_0_source1_matchingTag_bits_w_id ? buffer_12_valueReady : _GEN_1597; // @[ReorderBuffer.scala 160:{35,35}]
  wire  _GEN_1599 = 4'hd == io_decoders_0_source1_matchingTag_bits_w_id ? buffer_13_valueReady : _GEN_1598; // @[ReorderBuffer.scala 160:{35,35}]
  wire  _GEN_1600 = 4'he == io_decoders_0_source1_matchingTag_bits_w_id ? buffer_14_valueReady : _GEN_1599; // @[ReorderBuffer.scala 160:{35,35}]
  wire  _GEN_1601 = 4'hf == io_decoders_0_source1_matchingTag_bits_w_id ? buffer_15_valueReady : _GEN_1600; // @[ReorderBuffer.scala 160:{35,35}]
  wire [63:0] _GEN_1603 = 4'h1 == io_decoders_0_source1_matchingTag_bits_w_id ? buffer_1_value : buffer_0_value; // @[ReorderBuffer.scala 161:{34,34}]
  wire [63:0] _GEN_1604 = 4'h2 == io_decoders_0_source1_matchingTag_bits_w_id ? buffer_2_value : _GEN_1603; // @[ReorderBuffer.scala 161:{34,34}]
  wire [63:0] _GEN_1605 = 4'h3 == io_decoders_0_source1_matchingTag_bits_w_id ? buffer_3_value : _GEN_1604; // @[ReorderBuffer.scala 161:{34,34}]
  wire [63:0] _GEN_1606 = 4'h4 == io_decoders_0_source1_matchingTag_bits_w_id ? buffer_4_value : _GEN_1605; // @[ReorderBuffer.scala 161:{34,34}]
  wire [63:0] _GEN_1607 = 4'h5 == io_decoders_0_source1_matchingTag_bits_w_id ? buffer_5_value : _GEN_1606; // @[ReorderBuffer.scala 161:{34,34}]
  wire [63:0] _GEN_1608 = 4'h6 == io_decoders_0_source1_matchingTag_bits_w_id ? buffer_6_value : _GEN_1607; // @[ReorderBuffer.scala 161:{34,34}]
  wire [63:0] _GEN_1609 = 4'h7 == io_decoders_0_source1_matchingTag_bits_w_id ? buffer_7_value : _GEN_1608; // @[ReorderBuffer.scala 161:{34,34}]
  wire [63:0] _GEN_1610 = 4'h8 == io_decoders_0_source1_matchingTag_bits_w_id ? buffer_8_value : _GEN_1609; // @[ReorderBuffer.scala 161:{34,34}]
  wire [63:0] _GEN_1611 = 4'h9 == io_decoders_0_source1_matchingTag_bits_w_id ? buffer_9_value : _GEN_1610; // @[ReorderBuffer.scala 161:{34,34}]
  wire [63:0] _GEN_1612 = 4'ha == io_decoders_0_source1_matchingTag_bits_w_id ? buffer_10_value : _GEN_1611; // @[ReorderBuffer.scala 161:{34,34}]
  wire [63:0] _GEN_1613 = 4'hb == io_decoders_0_source1_matchingTag_bits_w_id ? buffer_11_value : _GEN_1612; // @[ReorderBuffer.scala 161:{34,34}]
  wire [63:0] _GEN_1614 = 4'hc == io_decoders_0_source1_matchingTag_bits_w_id ? buffer_12_value : _GEN_1613; // @[ReorderBuffer.scala 161:{34,34}]
  wire [63:0] _GEN_1615 = 4'hd == io_decoders_0_source1_matchingTag_bits_w_id ? buffer_13_value : _GEN_1614; // @[ReorderBuffer.scala 161:{34,34}]
  wire [63:0] _GEN_1616 = 4'he == io_decoders_0_source1_matchingTag_bits_w_id ? buffer_14_value : _GEN_1615; // @[ReorderBuffer.scala 161:{34,34}]
  wire [63:0] _GEN_1617 = 4'hf == io_decoders_0_source1_matchingTag_bits_w_id ? buffer_15_value : _GEN_1616; // @[ReorderBuffer.scala 161:{34,34}]
  wire  _GEN_1625 = 5'h2 == io_decoders_0_source2_sourceRegister ? registerTagMap_2_valid : 5'h1 ==
    io_decoders_0_source2_sourceRegister & registerTagMap_1_valid; // @[ReorderBuffer.scala 172:{41,41}]
  wire  _GEN_1626 = 5'h3 == io_decoders_0_source2_sourceRegister ? registerTagMap_3_valid : _GEN_1625; // @[ReorderBuffer.scala 172:{41,41}]
  wire  _GEN_1627 = 5'h4 == io_decoders_0_source2_sourceRegister ? registerTagMap_4_valid : _GEN_1626; // @[ReorderBuffer.scala 172:{41,41}]
  wire  _GEN_1628 = 5'h5 == io_decoders_0_source2_sourceRegister ? registerTagMap_5_valid : _GEN_1627; // @[ReorderBuffer.scala 172:{41,41}]
  wire  _GEN_1629 = 5'h6 == io_decoders_0_source2_sourceRegister ? registerTagMap_6_valid : _GEN_1628; // @[ReorderBuffer.scala 172:{41,41}]
  wire  _GEN_1630 = 5'h7 == io_decoders_0_source2_sourceRegister ? registerTagMap_7_valid : _GEN_1629; // @[ReorderBuffer.scala 172:{41,41}]
  wire  _GEN_1631 = 5'h8 == io_decoders_0_source2_sourceRegister ? registerTagMap_8_valid : _GEN_1630; // @[ReorderBuffer.scala 172:{41,41}]
  wire  _GEN_1632 = 5'h9 == io_decoders_0_source2_sourceRegister ? registerTagMap_9_valid : _GEN_1631; // @[ReorderBuffer.scala 172:{41,41}]
  wire  _GEN_1633 = 5'ha == io_decoders_0_source2_sourceRegister ? registerTagMap_10_valid : _GEN_1632; // @[ReorderBuffer.scala 172:{41,41}]
  wire  _GEN_1634 = 5'hb == io_decoders_0_source2_sourceRegister ? registerTagMap_11_valid : _GEN_1633; // @[ReorderBuffer.scala 172:{41,41}]
  wire  _GEN_1635 = 5'hc == io_decoders_0_source2_sourceRegister ? registerTagMap_12_valid : _GEN_1634; // @[ReorderBuffer.scala 172:{41,41}]
  wire  _GEN_1636 = 5'hd == io_decoders_0_source2_sourceRegister ? registerTagMap_13_valid : _GEN_1635; // @[ReorderBuffer.scala 172:{41,41}]
  wire  _GEN_1637 = 5'he == io_decoders_0_source2_sourceRegister ? registerTagMap_14_valid : _GEN_1636; // @[ReorderBuffer.scala 172:{41,41}]
  wire  _GEN_1638 = 5'hf == io_decoders_0_source2_sourceRegister ? registerTagMap_15_valid : _GEN_1637; // @[ReorderBuffer.scala 172:{41,41}]
  wire  _GEN_1639 = 5'h10 == io_decoders_0_source2_sourceRegister ? registerTagMap_16_valid : _GEN_1638; // @[ReorderBuffer.scala 172:{41,41}]
  wire  _GEN_1640 = 5'h11 == io_decoders_0_source2_sourceRegister ? registerTagMap_17_valid : _GEN_1639; // @[ReorderBuffer.scala 172:{41,41}]
  wire  _GEN_1641 = 5'h12 == io_decoders_0_source2_sourceRegister ? registerTagMap_18_valid : _GEN_1640; // @[ReorderBuffer.scala 172:{41,41}]
  wire  _GEN_1642 = 5'h13 == io_decoders_0_source2_sourceRegister ? registerTagMap_19_valid : _GEN_1641; // @[ReorderBuffer.scala 172:{41,41}]
  wire  _GEN_1643 = 5'h14 == io_decoders_0_source2_sourceRegister ? registerTagMap_20_valid : _GEN_1642; // @[ReorderBuffer.scala 172:{41,41}]
  wire  _GEN_1644 = 5'h15 == io_decoders_0_source2_sourceRegister ? registerTagMap_21_valid : _GEN_1643; // @[ReorderBuffer.scala 172:{41,41}]
  wire  _GEN_1645 = 5'h16 == io_decoders_0_source2_sourceRegister ? registerTagMap_22_valid : _GEN_1644; // @[ReorderBuffer.scala 172:{41,41}]
  wire  _GEN_1646 = 5'h17 == io_decoders_0_source2_sourceRegister ? registerTagMap_23_valid : _GEN_1645; // @[ReorderBuffer.scala 172:{41,41}]
  wire  _GEN_1647 = 5'h18 == io_decoders_0_source2_sourceRegister ? registerTagMap_24_valid : _GEN_1646; // @[ReorderBuffer.scala 172:{41,41}]
  wire  _GEN_1648 = 5'h19 == io_decoders_0_source2_sourceRegister ? registerTagMap_25_valid : _GEN_1647; // @[ReorderBuffer.scala 172:{41,41}]
  wire  _GEN_1649 = 5'h1a == io_decoders_0_source2_sourceRegister ? registerTagMap_26_valid : _GEN_1648; // @[ReorderBuffer.scala 172:{41,41}]
  wire  _GEN_1650 = 5'h1b == io_decoders_0_source2_sourceRegister ? registerTagMap_27_valid : _GEN_1649; // @[ReorderBuffer.scala 172:{41,41}]
  wire  _GEN_1651 = 5'h1c == io_decoders_0_source2_sourceRegister ? registerTagMap_28_valid : _GEN_1650; // @[ReorderBuffer.scala 172:{41,41}]
  wire  _GEN_1652 = 5'h1d == io_decoders_0_source2_sourceRegister ? registerTagMap_29_valid : _GEN_1651; // @[ReorderBuffer.scala 172:{41,41}]
  wire  _GEN_1653 = 5'h1e == io_decoders_0_source2_sourceRegister ? registerTagMap_30_valid : _GEN_1652; // @[ReorderBuffer.scala 172:{41,41}]
  wire  _GEN_1654 = 5'h1f == io_decoders_0_source2_sourceRegister ? registerTagMap_31_valid : _GEN_1653; // @[ReorderBuffer.scala 172:{41,41}]
  wire [3:0] _GEN_1656 = 5'h1 == io_decoders_0_source2_sourceRegister ? registerTagMap_1_tagId : 4'h0; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1657 = 5'h2 == io_decoders_0_source2_sourceRegister ? registerTagMap_2_tagId : _GEN_1656; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1658 = 5'h3 == io_decoders_0_source2_sourceRegister ? registerTagMap_3_tagId : _GEN_1657; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1659 = 5'h4 == io_decoders_0_source2_sourceRegister ? registerTagMap_4_tagId : _GEN_1658; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1660 = 5'h5 == io_decoders_0_source2_sourceRegister ? registerTagMap_5_tagId : _GEN_1659; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1661 = 5'h6 == io_decoders_0_source2_sourceRegister ? registerTagMap_6_tagId : _GEN_1660; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1662 = 5'h7 == io_decoders_0_source2_sourceRegister ? registerTagMap_7_tagId : _GEN_1661; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1663 = 5'h8 == io_decoders_0_source2_sourceRegister ? registerTagMap_8_tagId : _GEN_1662; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1664 = 5'h9 == io_decoders_0_source2_sourceRegister ? registerTagMap_9_tagId : _GEN_1663; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1665 = 5'ha == io_decoders_0_source2_sourceRegister ? registerTagMap_10_tagId : _GEN_1664; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1666 = 5'hb == io_decoders_0_source2_sourceRegister ? registerTagMap_11_tagId : _GEN_1665; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1667 = 5'hc == io_decoders_0_source2_sourceRegister ? registerTagMap_12_tagId : _GEN_1666; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1668 = 5'hd == io_decoders_0_source2_sourceRegister ? registerTagMap_13_tagId : _GEN_1667; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1669 = 5'he == io_decoders_0_source2_sourceRegister ? registerTagMap_14_tagId : _GEN_1668; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1670 = 5'hf == io_decoders_0_source2_sourceRegister ? registerTagMap_15_tagId : _GEN_1669; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1671 = 5'h10 == io_decoders_0_source2_sourceRegister ? registerTagMap_16_tagId : _GEN_1670; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1672 = 5'h11 == io_decoders_0_source2_sourceRegister ? registerTagMap_17_tagId : _GEN_1671; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1673 = 5'h12 == io_decoders_0_source2_sourceRegister ? registerTagMap_18_tagId : _GEN_1672; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1674 = 5'h13 == io_decoders_0_source2_sourceRegister ? registerTagMap_19_tagId : _GEN_1673; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1675 = 5'h14 == io_decoders_0_source2_sourceRegister ? registerTagMap_20_tagId : _GEN_1674; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1676 = 5'h15 == io_decoders_0_source2_sourceRegister ? registerTagMap_21_tagId : _GEN_1675; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1677 = 5'h16 == io_decoders_0_source2_sourceRegister ? registerTagMap_22_tagId : _GEN_1676; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1678 = 5'h17 == io_decoders_0_source2_sourceRegister ? registerTagMap_23_tagId : _GEN_1677; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1679 = 5'h18 == io_decoders_0_source2_sourceRegister ? registerTagMap_24_tagId : _GEN_1678; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1680 = 5'h19 == io_decoders_0_source2_sourceRegister ? registerTagMap_25_tagId : _GEN_1679; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1681 = 5'h1a == io_decoders_0_source2_sourceRegister ? registerTagMap_26_tagId : _GEN_1680; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1682 = 5'h1b == io_decoders_0_source2_sourceRegister ? registerTagMap_27_tagId : _GEN_1681; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1683 = 5'h1c == io_decoders_0_source2_sourceRegister ? registerTagMap_28_tagId : _GEN_1682; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1684 = 5'h1d == io_decoders_0_source2_sourceRegister ? registerTagMap_29_tagId : _GEN_1683; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1685 = 5'h1e == io_decoders_0_source2_sourceRegister ? registerTagMap_30_tagId : _GEN_1684; // @[Tag.scala 23:{10,10}]
  wire [3:0] io_decoders_0_source2_matchingTag_bits_w_id = 5'h1f == io_decoders_0_source2_sourceRegister ?
    registerTagMap_31_tagId : _GEN_1685; // @[Tag.scala 23:{10,10}]
  wire  _GEN_1688 = 4'h1 == io_decoders_0_source2_matchingTag_bits_w_id ? buffer_1_valueReady : buffer_0_valueReady; // @[ReorderBuffer.scala 177:{35,35}]
  wire  _GEN_1689 = 4'h2 == io_decoders_0_source2_matchingTag_bits_w_id ? buffer_2_valueReady : _GEN_1688; // @[ReorderBuffer.scala 177:{35,35}]
  wire  _GEN_1690 = 4'h3 == io_decoders_0_source2_matchingTag_bits_w_id ? buffer_3_valueReady : _GEN_1689; // @[ReorderBuffer.scala 177:{35,35}]
  wire  _GEN_1691 = 4'h4 == io_decoders_0_source2_matchingTag_bits_w_id ? buffer_4_valueReady : _GEN_1690; // @[ReorderBuffer.scala 177:{35,35}]
  wire  _GEN_1692 = 4'h5 == io_decoders_0_source2_matchingTag_bits_w_id ? buffer_5_valueReady : _GEN_1691; // @[ReorderBuffer.scala 177:{35,35}]
  wire  _GEN_1693 = 4'h6 == io_decoders_0_source2_matchingTag_bits_w_id ? buffer_6_valueReady : _GEN_1692; // @[ReorderBuffer.scala 177:{35,35}]
  wire  _GEN_1694 = 4'h7 == io_decoders_0_source2_matchingTag_bits_w_id ? buffer_7_valueReady : _GEN_1693; // @[ReorderBuffer.scala 177:{35,35}]
  wire  _GEN_1695 = 4'h8 == io_decoders_0_source2_matchingTag_bits_w_id ? buffer_8_valueReady : _GEN_1694; // @[ReorderBuffer.scala 177:{35,35}]
  wire  _GEN_1696 = 4'h9 == io_decoders_0_source2_matchingTag_bits_w_id ? buffer_9_valueReady : _GEN_1695; // @[ReorderBuffer.scala 177:{35,35}]
  wire  _GEN_1697 = 4'ha == io_decoders_0_source2_matchingTag_bits_w_id ? buffer_10_valueReady : _GEN_1696; // @[ReorderBuffer.scala 177:{35,35}]
  wire  _GEN_1698 = 4'hb == io_decoders_0_source2_matchingTag_bits_w_id ? buffer_11_valueReady : _GEN_1697; // @[ReorderBuffer.scala 177:{35,35}]
  wire  _GEN_1699 = 4'hc == io_decoders_0_source2_matchingTag_bits_w_id ? buffer_12_valueReady : _GEN_1698; // @[ReorderBuffer.scala 177:{35,35}]
  wire  _GEN_1700 = 4'hd == io_decoders_0_source2_matchingTag_bits_w_id ? buffer_13_valueReady : _GEN_1699; // @[ReorderBuffer.scala 177:{35,35}]
  wire  _GEN_1701 = 4'he == io_decoders_0_source2_matchingTag_bits_w_id ? buffer_14_valueReady : _GEN_1700; // @[ReorderBuffer.scala 177:{35,35}]
  wire  _GEN_1702 = 4'hf == io_decoders_0_source2_matchingTag_bits_w_id ? buffer_15_valueReady : _GEN_1701; // @[ReorderBuffer.scala 177:{35,35}]
  wire [63:0] _GEN_1704 = 4'h1 == io_decoders_0_source2_matchingTag_bits_w_id ? buffer_1_value : buffer_0_value; // @[ReorderBuffer.scala 178:{34,34}]
  wire [63:0] _GEN_1705 = 4'h2 == io_decoders_0_source2_matchingTag_bits_w_id ? buffer_2_value : _GEN_1704; // @[ReorderBuffer.scala 178:{34,34}]
  wire [63:0] _GEN_1706 = 4'h3 == io_decoders_0_source2_matchingTag_bits_w_id ? buffer_3_value : _GEN_1705; // @[ReorderBuffer.scala 178:{34,34}]
  wire [63:0] _GEN_1707 = 4'h4 == io_decoders_0_source2_matchingTag_bits_w_id ? buffer_4_value : _GEN_1706; // @[ReorderBuffer.scala 178:{34,34}]
  wire [63:0] _GEN_1708 = 4'h5 == io_decoders_0_source2_matchingTag_bits_w_id ? buffer_5_value : _GEN_1707; // @[ReorderBuffer.scala 178:{34,34}]
  wire [63:0] _GEN_1709 = 4'h6 == io_decoders_0_source2_matchingTag_bits_w_id ? buffer_6_value : _GEN_1708; // @[ReorderBuffer.scala 178:{34,34}]
  wire [63:0] _GEN_1710 = 4'h7 == io_decoders_0_source2_matchingTag_bits_w_id ? buffer_7_value : _GEN_1709; // @[ReorderBuffer.scala 178:{34,34}]
  wire [63:0] _GEN_1711 = 4'h8 == io_decoders_0_source2_matchingTag_bits_w_id ? buffer_8_value : _GEN_1710; // @[ReorderBuffer.scala 178:{34,34}]
  wire [63:0] _GEN_1712 = 4'h9 == io_decoders_0_source2_matchingTag_bits_w_id ? buffer_9_value : _GEN_1711; // @[ReorderBuffer.scala 178:{34,34}]
  wire [63:0] _GEN_1713 = 4'ha == io_decoders_0_source2_matchingTag_bits_w_id ? buffer_10_value : _GEN_1712; // @[ReorderBuffer.scala 178:{34,34}]
  wire [63:0] _GEN_1714 = 4'hb == io_decoders_0_source2_matchingTag_bits_w_id ? buffer_11_value : _GEN_1713; // @[ReorderBuffer.scala 178:{34,34}]
  wire [63:0] _GEN_1715 = 4'hc == io_decoders_0_source2_matchingTag_bits_w_id ? buffer_12_value : _GEN_1714; // @[ReorderBuffer.scala 178:{34,34}]
  wire [63:0] _GEN_1716 = 4'hd == io_decoders_0_source2_matchingTag_bits_w_id ? buffer_13_value : _GEN_1715; // @[ReorderBuffer.scala 178:{34,34}]
  wire [63:0] _GEN_1717 = 4'he == io_decoders_0_source2_matchingTag_bits_w_id ? buffer_14_value : _GEN_1716; // @[ReorderBuffer.scala 178:{34,34}]
  wire [63:0] _GEN_1718 = 4'hf == io_decoders_0_source2_matchingTag_bits_w_id ? buffer_15_value : _GEN_1717; // @[ReorderBuffer.scala 178:{34,34}]
  wire [3:0] _GEN_1853 = {{1'd0}, tailDelta}; // @[ReorderBuffer.scala 193:45]
  wire [3:0] _tail_T_1 = tail + _GEN_1853; // @[ReorderBuffer.scala 193:45]
  wire [2:0] _io_csr_retireCount_T = io_isError ? 3'h0 : tailDelta; // @[ReorderBuffer.scala 194:28]
  wire  _T_19 = io_collectedOutputs_outputs_valid & ~io_collectedOutputs_outputs_bits_resultType & ~
    io_collectedOutputs_outputs_bits_tag_threadId; // @[ReorderBuffer.scala 200:68]
  wire  _GEN_1756 = 4'h0 == io_collectedOutputs_outputs_bits_tag_id | _GEN_1314; // @[ReorderBuffer.scala 204:{43,43}]
  wire  _GEN_1757 = 4'h1 == io_collectedOutputs_outputs_bits_tag_id | _GEN_1315; // @[ReorderBuffer.scala 204:{43,43}]
  wire  _GEN_1758 = 4'h2 == io_collectedOutputs_outputs_bits_tag_id | _GEN_1316; // @[ReorderBuffer.scala 204:{43,43}]
  wire  _GEN_1759 = 4'h3 == io_collectedOutputs_outputs_bits_tag_id | _GEN_1317; // @[ReorderBuffer.scala 204:{43,43}]
  wire  _GEN_1760 = 4'h4 == io_collectedOutputs_outputs_bits_tag_id | _GEN_1318; // @[ReorderBuffer.scala 204:{43,43}]
  wire  _GEN_1761 = 4'h5 == io_collectedOutputs_outputs_bits_tag_id | _GEN_1319; // @[ReorderBuffer.scala 204:{43,43}]
  wire  _GEN_1762 = 4'h6 == io_collectedOutputs_outputs_bits_tag_id | _GEN_1320; // @[ReorderBuffer.scala 204:{43,43}]
  wire  _GEN_1763 = 4'h7 == io_collectedOutputs_outputs_bits_tag_id | _GEN_1321; // @[ReorderBuffer.scala 204:{43,43}]
  wire  _GEN_1764 = 4'h8 == io_collectedOutputs_outputs_bits_tag_id | _GEN_1322; // @[ReorderBuffer.scala 204:{43,43}]
  wire  _GEN_1765 = 4'h9 == io_collectedOutputs_outputs_bits_tag_id | _GEN_1323; // @[ReorderBuffer.scala 204:{43,43}]
  wire  _GEN_1766 = 4'ha == io_collectedOutputs_outputs_bits_tag_id | _GEN_1324; // @[ReorderBuffer.scala 204:{43,43}]
  wire  _GEN_1767 = 4'hb == io_collectedOutputs_outputs_bits_tag_id | _GEN_1325; // @[ReorderBuffer.scala 204:{43,43}]
  wire  _GEN_1768 = 4'hc == io_collectedOutputs_outputs_bits_tag_id | _GEN_1326; // @[ReorderBuffer.scala 204:{43,43}]
  wire  _GEN_1769 = 4'hd == io_collectedOutputs_outputs_bits_tag_id | _GEN_1327; // @[ReorderBuffer.scala 204:{43,43}]
  wire  _GEN_1770 = 4'he == io_collectedOutputs_outputs_bits_tag_id | _GEN_1328; // @[ReorderBuffer.scala 204:{43,43}]
  wire  _GEN_1771 = 4'hf == io_collectedOutputs_outputs_bits_tag_id | _GEN_1329; // @[ReorderBuffer.scala 204:{43,43}]
  assign io_decoders_0_source1_matchingTag_valid = io_decoders_0_source1_sourceRegister != 5'h0 & _GEN_1553; // @[ReorderBuffer.scala 151:50 155:41 163:41]
  assign io_decoders_0_source1_matchingTag_bits_id = io_decoders_0_source1_sourceRegister != 5'h0 ?
    io_decoders_0_source1_matchingTag_bits_w_id : 4'h0; // @[ReorderBuffer.scala 151:50 156:40 164:40]
  assign io_decoders_0_source1_value_valid = io_decoders_0_source1_sourceRegister != 5'h0 & _GEN_1601; // @[ReorderBuffer.scala 151:50 160:35 165:35]
  assign io_decoders_0_source1_value_bits = io_decoders_0_source1_sourceRegister != 5'h0 ? _GEN_1617 : 64'h0; // @[ReorderBuffer.scala 151:50 161:34 166:34]
  assign io_decoders_0_source2_matchingTag_valid = io_decoders_0_source2_sourceRegister != 5'h0 & _GEN_1654; // @[ReorderBuffer.scala 169:50 172:41 180:41]
  assign io_decoders_0_source2_matchingTag_bits_id = io_decoders_0_source2_sourceRegister != 5'h0 ?
    io_decoders_0_source2_matchingTag_bits_w_id : 4'h0; // @[ReorderBuffer.scala 169:50 173:40 181:40]
  assign io_decoders_0_source2_value_valid = io_decoders_0_source2_sourceRegister != 5'h0 & _GEN_1702; // @[ReorderBuffer.scala 169:50 177:35 182:35]
  assign io_decoders_0_source2_value_bits = io_decoders_0_source2_sourceRegister != 5'h0 ? _GEN_1718 : 64'h0; // @[ReorderBuffer.scala 169:50 178:34 183:34]
  assign io_decoders_0_destination_destinationTag_id = head; // @[Tag.scala 21:17 23:10]
  assign io_decoders_0_ready = _io_decoders_0_ready_T_1 != tail; // @[ReorderBuffer.scala 129:55]
  assign io_registerFile_0_valid = canCommit & ~_GEN_47; // @[ReorderBuffer.scala 83:27]
  assign io_registerFile_0_bits_destinationRegister = canCommit ? _GEN_209 : 5'h0; // @[ReorderBuffer.scala 88:21 85:33]
  assign io_registerFile_0_bits_value = canCommit ? _GEN_208 : 64'h0; // @[ReorderBuffer.scala 84:19 88:21]
  assign io_registerFile_1_valid = canCommit_1 & ~_GEN_346; // @[ReorderBuffer.scala 83:27]
  assign io_registerFile_1_bits_destinationRegister = canCommit_1 ? _GEN_508 : 5'h0; // @[ReorderBuffer.scala 88:21 85:33]
  assign io_registerFile_1_bits_value = canCommit_1 ? _GEN_507 : 64'h0; // @[ReorderBuffer.scala 84:19 88:21]
  assign io_registerFile_2_valid = canCommit_2 & ~_GEN_647; // @[ReorderBuffer.scala 83:27]
  assign io_registerFile_2_bits_destinationRegister = canCommit_2 ? _GEN_809 : 5'h0; // @[ReorderBuffer.scala 88:21 85:33]
  assign io_registerFile_2_bits_value = canCommit_2 ? _GEN_808 : 64'h0; // @[ReorderBuffer.scala 84:19 88:21]
  assign io_registerFile_3_valid = canCommit_3 & ~_GEN_948; // @[ReorderBuffer.scala 83:27]
  assign io_registerFile_3_bits_destinationRegister = canCommit_3 ? _GEN_1110 : 5'h0; // @[ReorderBuffer.scala 88:21 85:33]
  assign io_registerFile_3_bits_value = canCommit_3 ? _GEN_1109 : 64'h0; // @[ReorderBuffer.scala 84:19 88:21]
  assign io_loadStoreQueue_0_valid = canCommit & _GEN_31; // @[ReorderBuffer.scala 106:21 109:17 113:17]
  assign io_loadStoreQueue_0_bits_destinationTag_id = canCommit ? index : 4'h0; // @[ReorderBuffer.scala 106:21 108:31 112:31]
  assign io_loadStoreQueue_1_valid = canCommit_1 & _GEN_330; // @[ReorderBuffer.scala 106:21 109:17 113:17]
  assign io_loadStoreQueue_1_bits_destinationTag_id = canCommit_1 ? index_1 : 4'h0; // @[ReorderBuffer.scala 106:21 108:31 112:31]
  assign io_loadStoreQueue_2_valid = canCommit_2 & _GEN_631; // @[ReorderBuffer.scala 106:21 109:17 113:17]
  assign io_loadStoreQueue_2_bits_destinationTag_id = canCommit_2 ? index_2 : 4'h0; // @[ReorderBuffer.scala 106:21 108:31 112:31]
  assign io_loadStoreQueue_3_valid = canCommit_3 & _GEN_932; // @[ReorderBuffer.scala 106:21 109:17 113:17]
  assign io_loadStoreQueue_3_bits_destinationTag_id = canCommit_3 ? index_3 : 4'h0; // @[ReorderBuffer.scala 106:21 108:31 112:31]
  assign io_isEmpty = head == tail; // @[ReorderBuffer.scala 195:22]
  assign io_csr_retireCount = _io_csr_retireCount_T[1:0]; // @[ReorderBuffer.scala 194:22]
  assign io_isError = canCommit_3 ? _GEN_1145 : _GEN_881; // @[ReorderBuffer.scala 88:21]
  always @(posedge clock) begin
    if (reset) begin // @[ReorderBuffer.scala 53:21]
      head <= 4'h0; // @[ReorderBuffer.scala 53:21]
    end else if (_T_8) begin // @[ReorderBuffer.scala 189:10]
      head <= _io_decoders_0_ready_T_1;
    end
    if (reset) begin // @[ReorderBuffer.scala 54:21]
      tail <= 4'h0; // @[ReorderBuffer.scala 54:21]
    end else if (io_isError) begin // @[ReorderBuffer.scala 193:14]
      if (_T_8) begin // @[ReorderBuffer.scala 189:10]
        tail <= _io_decoders_0_ready_T_1;
      end else begin
        tail <= head;
      end
    end else begin
      tail <= _tail_T_1;
    end
    if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'h0 == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_0_destinationRegister <= io_decoders_0_destination_destinationRegister; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      buffer_0_valueReady <= _GEN_1756;
    end else if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'h0 == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_0_valueReady <= 1'h0; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      if (4'h0 == io_collectedOutputs_outputs_bits_tag_id) begin // @[ReorderBuffer.scala 202:38]
        buffer_0_value <= io_collectedOutputs_outputs_bits_value; // @[ReorderBuffer.scala 202:38]
      end else begin
        buffer_0_value <= _GEN_1330;
      end
    end else begin
      buffer_0_value <= _GEN_1330;
    end
    if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'h0 == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_0_storeSign <= io_decoders_0_destination_storeSign; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      if (4'h0 == io_collectedOutputs_outputs_bits_tag_id) begin // @[ReorderBuffer.scala 203:40]
        buffer_0_isError <= io_collectedOutputs_outputs_bits_isError; // @[ReorderBuffer.scala 203:40]
      end else begin
        buffer_0_isError <= _GEN_1378;
      end
    end else begin
      buffer_0_isError <= _GEN_1378;
    end
    if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'h1 == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_1_destinationRegister <= io_decoders_0_destination_destinationRegister; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      buffer_1_valueReady <= _GEN_1757;
    end else if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'h1 == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_1_valueReady <= 1'h0; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      if (4'h1 == io_collectedOutputs_outputs_bits_tag_id) begin // @[ReorderBuffer.scala 202:38]
        buffer_1_value <= io_collectedOutputs_outputs_bits_value; // @[ReorderBuffer.scala 202:38]
      end else begin
        buffer_1_value <= _GEN_1331;
      end
    end else begin
      buffer_1_value <= _GEN_1331;
    end
    if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'h1 == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_1_storeSign <= io_decoders_0_destination_storeSign; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      if (4'h1 == io_collectedOutputs_outputs_bits_tag_id) begin // @[ReorderBuffer.scala 203:40]
        buffer_1_isError <= io_collectedOutputs_outputs_bits_isError; // @[ReorderBuffer.scala 203:40]
      end else begin
        buffer_1_isError <= _GEN_1379;
      end
    end else begin
      buffer_1_isError <= _GEN_1379;
    end
    if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'h2 == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_2_destinationRegister <= io_decoders_0_destination_destinationRegister; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      buffer_2_valueReady <= _GEN_1758;
    end else if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'h2 == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_2_valueReady <= 1'h0; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      if (4'h2 == io_collectedOutputs_outputs_bits_tag_id) begin // @[ReorderBuffer.scala 202:38]
        buffer_2_value <= io_collectedOutputs_outputs_bits_value; // @[ReorderBuffer.scala 202:38]
      end else begin
        buffer_2_value <= _GEN_1332;
      end
    end else begin
      buffer_2_value <= _GEN_1332;
    end
    if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'h2 == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_2_storeSign <= io_decoders_0_destination_storeSign; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      if (4'h2 == io_collectedOutputs_outputs_bits_tag_id) begin // @[ReorderBuffer.scala 203:40]
        buffer_2_isError <= io_collectedOutputs_outputs_bits_isError; // @[ReorderBuffer.scala 203:40]
      end else begin
        buffer_2_isError <= _GEN_1380;
      end
    end else begin
      buffer_2_isError <= _GEN_1380;
    end
    if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'h3 == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_3_destinationRegister <= io_decoders_0_destination_destinationRegister; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      buffer_3_valueReady <= _GEN_1759;
    end else if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'h3 == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_3_valueReady <= 1'h0; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      if (4'h3 == io_collectedOutputs_outputs_bits_tag_id) begin // @[ReorderBuffer.scala 202:38]
        buffer_3_value <= io_collectedOutputs_outputs_bits_value; // @[ReorderBuffer.scala 202:38]
      end else begin
        buffer_3_value <= _GEN_1333;
      end
    end else begin
      buffer_3_value <= _GEN_1333;
    end
    if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'h3 == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_3_storeSign <= io_decoders_0_destination_storeSign; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      if (4'h3 == io_collectedOutputs_outputs_bits_tag_id) begin // @[ReorderBuffer.scala 203:40]
        buffer_3_isError <= io_collectedOutputs_outputs_bits_isError; // @[ReorderBuffer.scala 203:40]
      end else begin
        buffer_3_isError <= _GEN_1381;
      end
    end else begin
      buffer_3_isError <= _GEN_1381;
    end
    if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'h4 == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_4_destinationRegister <= io_decoders_0_destination_destinationRegister; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      buffer_4_valueReady <= _GEN_1760;
    end else if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'h4 == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_4_valueReady <= 1'h0; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      if (4'h4 == io_collectedOutputs_outputs_bits_tag_id) begin // @[ReorderBuffer.scala 202:38]
        buffer_4_value <= io_collectedOutputs_outputs_bits_value; // @[ReorderBuffer.scala 202:38]
      end else begin
        buffer_4_value <= _GEN_1334;
      end
    end else begin
      buffer_4_value <= _GEN_1334;
    end
    if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'h4 == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_4_storeSign <= io_decoders_0_destination_storeSign; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      if (4'h4 == io_collectedOutputs_outputs_bits_tag_id) begin // @[ReorderBuffer.scala 203:40]
        buffer_4_isError <= io_collectedOutputs_outputs_bits_isError; // @[ReorderBuffer.scala 203:40]
      end else begin
        buffer_4_isError <= _GEN_1382;
      end
    end else begin
      buffer_4_isError <= _GEN_1382;
    end
    if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'h5 == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_5_destinationRegister <= io_decoders_0_destination_destinationRegister; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      buffer_5_valueReady <= _GEN_1761;
    end else if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'h5 == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_5_valueReady <= 1'h0; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      if (4'h5 == io_collectedOutputs_outputs_bits_tag_id) begin // @[ReorderBuffer.scala 202:38]
        buffer_5_value <= io_collectedOutputs_outputs_bits_value; // @[ReorderBuffer.scala 202:38]
      end else begin
        buffer_5_value <= _GEN_1335;
      end
    end else begin
      buffer_5_value <= _GEN_1335;
    end
    if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'h5 == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_5_storeSign <= io_decoders_0_destination_storeSign; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      if (4'h5 == io_collectedOutputs_outputs_bits_tag_id) begin // @[ReorderBuffer.scala 203:40]
        buffer_5_isError <= io_collectedOutputs_outputs_bits_isError; // @[ReorderBuffer.scala 203:40]
      end else begin
        buffer_5_isError <= _GEN_1383;
      end
    end else begin
      buffer_5_isError <= _GEN_1383;
    end
    if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'h6 == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_6_destinationRegister <= io_decoders_0_destination_destinationRegister; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      buffer_6_valueReady <= _GEN_1762;
    end else if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'h6 == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_6_valueReady <= 1'h0; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      if (4'h6 == io_collectedOutputs_outputs_bits_tag_id) begin // @[ReorderBuffer.scala 202:38]
        buffer_6_value <= io_collectedOutputs_outputs_bits_value; // @[ReorderBuffer.scala 202:38]
      end else begin
        buffer_6_value <= _GEN_1336;
      end
    end else begin
      buffer_6_value <= _GEN_1336;
    end
    if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'h6 == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_6_storeSign <= io_decoders_0_destination_storeSign; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      if (4'h6 == io_collectedOutputs_outputs_bits_tag_id) begin // @[ReorderBuffer.scala 203:40]
        buffer_6_isError <= io_collectedOutputs_outputs_bits_isError; // @[ReorderBuffer.scala 203:40]
      end else begin
        buffer_6_isError <= _GEN_1384;
      end
    end else begin
      buffer_6_isError <= _GEN_1384;
    end
    if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'h7 == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_7_destinationRegister <= io_decoders_0_destination_destinationRegister; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      buffer_7_valueReady <= _GEN_1763;
    end else if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'h7 == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_7_valueReady <= 1'h0; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      if (4'h7 == io_collectedOutputs_outputs_bits_tag_id) begin // @[ReorderBuffer.scala 202:38]
        buffer_7_value <= io_collectedOutputs_outputs_bits_value; // @[ReorderBuffer.scala 202:38]
      end else begin
        buffer_7_value <= _GEN_1337;
      end
    end else begin
      buffer_7_value <= _GEN_1337;
    end
    if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'h7 == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_7_storeSign <= io_decoders_0_destination_storeSign; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      if (4'h7 == io_collectedOutputs_outputs_bits_tag_id) begin // @[ReorderBuffer.scala 203:40]
        buffer_7_isError <= io_collectedOutputs_outputs_bits_isError; // @[ReorderBuffer.scala 203:40]
      end else begin
        buffer_7_isError <= _GEN_1385;
      end
    end else begin
      buffer_7_isError <= _GEN_1385;
    end
    if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'h8 == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_8_destinationRegister <= io_decoders_0_destination_destinationRegister; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      buffer_8_valueReady <= _GEN_1764;
    end else if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'h8 == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_8_valueReady <= 1'h0; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      if (4'h8 == io_collectedOutputs_outputs_bits_tag_id) begin // @[ReorderBuffer.scala 202:38]
        buffer_8_value <= io_collectedOutputs_outputs_bits_value; // @[ReorderBuffer.scala 202:38]
      end else begin
        buffer_8_value <= _GEN_1338;
      end
    end else begin
      buffer_8_value <= _GEN_1338;
    end
    if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'h8 == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_8_storeSign <= io_decoders_0_destination_storeSign; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      if (4'h8 == io_collectedOutputs_outputs_bits_tag_id) begin // @[ReorderBuffer.scala 203:40]
        buffer_8_isError <= io_collectedOutputs_outputs_bits_isError; // @[ReorderBuffer.scala 203:40]
      end else begin
        buffer_8_isError <= _GEN_1386;
      end
    end else begin
      buffer_8_isError <= _GEN_1386;
    end
    if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'h9 == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_9_destinationRegister <= io_decoders_0_destination_destinationRegister; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      buffer_9_valueReady <= _GEN_1765;
    end else if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'h9 == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_9_valueReady <= 1'h0; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      if (4'h9 == io_collectedOutputs_outputs_bits_tag_id) begin // @[ReorderBuffer.scala 202:38]
        buffer_9_value <= io_collectedOutputs_outputs_bits_value; // @[ReorderBuffer.scala 202:38]
      end else begin
        buffer_9_value <= _GEN_1339;
      end
    end else begin
      buffer_9_value <= _GEN_1339;
    end
    if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'h9 == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_9_storeSign <= io_decoders_0_destination_storeSign; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      if (4'h9 == io_collectedOutputs_outputs_bits_tag_id) begin // @[ReorderBuffer.scala 203:40]
        buffer_9_isError <= io_collectedOutputs_outputs_bits_isError; // @[ReorderBuffer.scala 203:40]
      end else begin
        buffer_9_isError <= _GEN_1387;
      end
    end else begin
      buffer_9_isError <= _GEN_1387;
    end
    if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'ha == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_10_destinationRegister <= io_decoders_0_destination_destinationRegister; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      buffer_10_valueReady <= _GEN_1766;
    end else if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'ha == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_10_valueReady <= 1'h0; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      if (4'ha == io_collectedOutputs_outputs_bits_tag_id) begin // @[ReorderBuffer.scala 202:38]
        buffer_10_value <= io_collectedOutputs_outputs_bits_value; // @[ReorderBuffer.scala 202:38]
      end else begin
        buffer_10_value <= _GEN_1340;
      end
    end else begin
      buffer_10_value <= _GEN_1340;
    end
    if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'ha == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_10_storeSign <= io_decoders_0_destination_storeSign; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      if (4'ha == io_collectedOutputs_outputs_bits_tag_id) begin // @[ReorderBuffer.scala 203:40]
        buffer_10_isError <= io_collectedOutputs_outputs_bits_isError; // @[ReorderBuffer.scala 203:40]
      end else begin
        buffer_10_isError <= _GEN_1388;
      end
    end else begin
      buffer_10_isError <= _GEN_1388;
    end
    if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'hb == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_11_destinationRegister <= io_decoders_0_destination_destinationRegister; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      buffer_11_valueReady <= _GEN_1767;
    end else if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'hb == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_11_valueReady <= 1'h0; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      if (4'hb == io_collectedOutputs_outputs_bits_tag_id) begin // @[ReorderBuffer.scala 202:38]
        buffer_11_value <= io_collectedOutputs_outputs_bits_value; // @[ReorderBuffer.scala 202:38]
      end else begin
        buffer_11_value <= _GEN_1341;
      end
    end else begin
      buffer_11_value <= _GEN_1341;
    end
    if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'hb == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_11_storeSign <= io_decoders_0_destination_storeSign; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      if (4'hb == io_collectedOutputs_outputs_bits_tag_id) begin // @[ReorderBuffer.scala 203:40]
        buffer_11_isError <= io_collectedOutputs_outputs_bits_isError; // @[ReorderBuffer.scala 203:40]
      end else begin
        buffer_11_isError <= _GEN_1389;
      end
    end else begin
      buffer_11_isError <= _GEN_1389;
    end
    if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'hc == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_12_destinationRegister <= io_decoders_0_destination_destinationRegister; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      buffer_12_valueReady <= _GEN_1768;
    end else if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'hc == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_12_valueReady <= 1'h0; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      if (4'hc == io_collectedOutputs_outputs_bits_tag_id) begin // @[ReorderBuffer.scala 202:38]
        buffer_12_value <= io_collectedOutputs_outputs_bits_value; // @[ReorderBuffer.scala 202:38]
      end else begin
        buffer_12_value <= _GEN_1342;
      end
    end else begin
      buffer_12_value <= _GEN_1342;
    end
    if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'hc == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_12_storeSign <= io_decoders_0_destination_storeSign; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      if (4'hc == io_collectedOutputs_outputs_bits_tag_id) begin // @[ReorderBuffer.scala 203:40]
        buffer_12_isError <= io_collectedOutputs_outputs_bits_isError; // @[ReorderBuffer.scala 203:40]
      end else begin
        buffer_12_isError <= _GEN_1390;
      end
    end else begin
      buffer_12_isError <= _GEN_1390;
    end
    if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'hd == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_13_destinationRegister <= io_decoders_0_destination_destinationRegister; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      buffer_13_valueReady <= _GEN_1769;
    end else if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'hd == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_13_valueReady <= 1'h0; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      if (4'hd == io_collectedOutputs_outputs_bits_tag_id) begin // @[ReorderBuffer.scala 202:38]
        buffer_13_value <= io_collectedOutputs_outputs_bits_value; // @[ReorderBuffer.scala 202:38]
      end else begin
        buffer_13_value <= _GEN_1343;
      end
    end else begin
      buffer_13_value <= _GEN_1343;
    end
    if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'hd == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_13_storeSign <= io_decoders_0_destination_storeSign; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      if (4'hd == io_collectedOutputs_outputs_bits_tag_id) begin // @[ReorderBuffer.scala 203:40]
        buffer_13_isError <= io_collectedOutputs_outputs_bits_isError; // @[ReorderBuffer.scala 203:40]
      end else begin
        buffer_13_isError <= _GEN_1391;
      end
    end else begin
      buffer_13_isError <= _GEN_1391;
    end
    if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'he == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_14_destinationRegister <= io_decoders_0_destination_destinationRegister; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      buffer_14_valueReady <= _GEN_1770;
    end else if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'he == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_14_valueReady <= 1'h0; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      if (4'he == io_collectedOutputs_outputs_bits_tag_id) begin // @[ReorderBuffer.scala 202:38]
        buffer_14_value <= io_collectedOutputs_outputs_bits_value; // @[ReorderBuffer.scala 202:38]
      end else begin
        buffer_14_value <= _GEN_1344;
      end
    end else begin
      buffer_14_value <= _GEN_1344;
    end
    if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'he == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_14_storeSign <= io_decoders_0_destination_storeSign; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      if (4'he == io_collectedOutputs_outputs_bits_tag_id) begin // @[ReorderBuffer.scala 203:40]
        buffer_14_isError <= io_collectedOutputs_outputs_bits_isError; // @[ReorderBuffer.scala 203:40]
      end else begin
        buffer_14_isError <= _GEN_1392;
      end
    end else begin
      buffer_14_isError <= _GEN_1392;
    end
    if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'hf == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_15_destinationRegister <= io_decoders_0_destination_destinationRegister; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      buffer_15_valueReady <= _GEN_1771;
    end else if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'hf == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_15_valueReady <= 1'h0; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      if (4'hf == io_collectedOutputs_outputs_bits_tag_id) begin // @[ReorderBuffer.scala 202:38]
        buffer_15_value <= io_collectedOutputs_outputs_bits_value; // @[ReorderBuffer.scala 202:38]
      end else begin
        buffer_15_value <= _GEN_1345;
      end
    end else begin
      buffer_15_value <= _GEN_1345;
    end
    if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'hf == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_15_storeSign <= io_decoders_0_destination_storeSign; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      if (4'hf == io_collectedOutputs_outputs_bits_tag_id) begin // @[ReorderBuffer.scala 203:40]
        buffer_15_isError <= io_collectedOutputs_outputs_bits_isError; // @[ReorderBuffer.scala 203:40]
      end else begin
        buffer_15_isError <= _GEN_1393;
      end
    end else begin
      buffer_15_isError <= _GEN_1393;
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_1_valid <= 1'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      registerTagMap_1_valid <= _GEN_1395;
    end else if (canCommit_3) begin // @[ReorderBuffer.scala 88:21]
      if (_io_registerFile_3_valid_T) begin // @[ReorderBuffer.scala 89:22]
        registerTagMap_1_valid <= _GEN_1078;
      end else begin
        registerTagMap_1_valid <= _GEN_848;
      end
    end else begin
      registerTagMap_1_valid <= _GEN_848;
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_1_tagId <= 4'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      if (5'h1 == io_decoders_0_destination_destinationRegister) begin // @[ReorderBuffer.scala 149:15]
        registerTagMap_1_tagId <= head; // @[ReorderBuffer.scala 149:15]
      end
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_2_valid <= 1'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      registerTagMap_2_valid <= _GEN_1396;
    end else if (canCommit_3) begin // @[ReorderBuffer.scala 88:21]
      if (_io_registerFile_3_valid_T) begin // @[ReorderBuffer.scala 89:22]
        registerTagMap_2_valid <= _GEN_1079;
      end else begin
        registerTagMap_2_valid <= _GEN_849;
      end
    end else begin
      registerTagMap_2_valid <= _GEN_849;
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_2_tagId <= 4'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      if (5'h2 == io_decoders_0_destination_destinationRegister) begin // @[ReorderBuffer.scala 149:15]
        registerTagMap_2_tagId <= head; // @[ReorderBuffer.scala 149:15]
      end
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_3_valid <= 1'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      registerTagMap_3_valid <= _GEN_1397;
    end else if (canCommit_3) begin // @[ReorderBuffer.scala 88:21]
      if (_io_registerFile_3_valid_T) begin // @[ReorderBuffer.scala 89:22]
        registerTagMap_3_valid <= _GEN_1080;
      end else begin
        registerTagMap_3_valid <= _GEN_850;
      end
    end else begin
      registerTagMap_3_valid <= _GEN_850;
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_3_tagId <= 4'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      if (5'h3 == io_decoders_0_destination_destinationRegister) begin // @[ReorderBuffer.scala 149:15]
        registerTagMap_3_tagId <= head; // @[ReorderBuffer.scala 149:15]
      end
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_4_valid <= 1'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      registerTagMap_4_valid <= _GEN_1398;
    end else if (canCommit_3) begin // @[ReorderBuffer.scala 88:21]
      if (_io_registerFile_3_valid_T) begin // @[ReorderBuffer.scala 89:22]
        registerTagMap_4_valid <= _GEN_1081;
      end else begin
        registerTagMap_4_valid <= _GEN_851;
      end
    end else begin
      registerTagMap_4_valid <= _GEN_851;
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_4_tagId <= 4'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      if (5'h4 == io_decoders_0_destination_destinationRegister) begin // @[ReorderBuffer.scala 149:15]
        registerTagMap_4_tagId <= head; // @[ReorderBuffer.scala 149:15]
      end
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_5_valid <= 1'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      registerTagMap_5_valid <= _GEN_1399;
    end else if (canCommit_3) begin // @[ReorderBuffer.scala 88:21]
      if (_io_registerFile_3_valid_T) begin // @[ReorderBuffer.scala 89:22]
        registerTagMap_5_valid <= _GEN_1082;
      end else begin
        registerTagMap_5_valid <= _GEN_852;
      end
    end else begin
      registerTagMap_5_valid <= _GEN_852;
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_5_tagId <= 4'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      if (5'h5 == io_decoders_0_destination_destinationRegister) begin // @[ReorderBuffer.scala 149:15]
        registerTagMap_5_tagId <= head; // @[ReorderBuffer.scala 149:15]
      end
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_6_valid <= 1'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      registerTagMap_6_valid <= _GEN_1400;
    end else if (canCommit_3) begin // @[ReorderBuffer.scala 88:21]
      if (_io_registerFile_3_valid_T) begin // @[ReorderBuffer.scala 89:22]
        registerTagMap_6_valid <= _GEN_1083;
      end else begin
        registerTagMap_6_valid <= _GEN_853;
      end
    end else begin
      registerTagMap_6_valid <= _GEN_853;
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_6_tagId <= 4'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      if (5'h6 == io_decoders_0_destination_destinationRegister) begin // @[ReorderBuffer.scala 149:15]
        registerTagMap_6_tagId <= head; // @[ReorderBuffer.scala 149:15]
      end
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_7_valid <= 1'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      registerTagMap_7_valid <= _GEN_1401;
    end else if (canCommit_3) begin // @[ReorderBuffer.scala 88:21]
      if (_io_registerFile_3_valid_T) begin // @[ReorderBuffer.scala 89:22]
        registerTagMap_7_valid <= _GEN_1084;
      end else begin
        registerTagMap_7_valid <= _GEN_854;
      end
    end else begin
      registerTagMap_7_valid <= _GEN_854;
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_7_tagId <= 4'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      if (5'h7 == io_decoders_0_destination_destinationRegister) begin // @[ReorderBuffer.scala 149:15]
        registerTagMap_7_tagId <= head; // @[ReorderBuffer.scala 149:15]
      end
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_8_valid <= 1'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      registerTagMap_8_valid <= _GEN_1402;
    end else if (canCommit_3) begin // @[ReorderBuffer.scala 88:21]
      if (_io_registerFile_3_valid_T) begin // @[ReorderBuffer.scala 89:22]
        registerTagMap_8_valid <= _GEN_1085;
      end else begin
        registerTagMap_8_valid <= _GEN_855;
      end
    end else begin
      registerTagMap_8_valid <= _GEN_855;
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_8_tagId <= 4'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      if (5'h8 == io_decoders_0_destination_destinationRegister) begin // @[ReorderBuffer.scala 149:15]
        registerTagMap_8_tagId <= head; // @[ReorderBuffer.scala 149:15]
      end
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_9_valid <= 1'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      registerTagMap_9_valid <= _GEN_1403;
    end else if (canCommit_3) begin // @[ReorderBuffer.scala 88:21]
      if (_io_registerFile_3_valid_T) begin // @[ReorderBuffer.scala 89:22]
        registerTagMap_9_valid <= _GEN_1086;
      end else begin
        registerTagMap_9_valid <= _GEN_856;
      end
    end else begin
      registerTagMap_9_valid <= _GEN_856;
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_9_tagId <= 4'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      if (5'h9 == io_decoders_0_destination_destinationRegister) begin // @[ReorderBuffer.scala 149:15]
        registerTagMap_9_tagId <= head; // @[ReorderBuffer.scala 149:15]
      end
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_10_valid <= 1'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      registerTagMap_10_valid <= _GEN_1404;
    end else if (canCommit_3) begin // @[ReorderBuffer.scala 88:21]
      if (_io_registerFile_3_valid_T) begin // @[ReorderBuffer.scala 89:22]
        registerTagMap_10_valid <= _GEN_1087;
      end else begin
        registerTagMap_10_valid <= _GEN_857;
      end
    end else begin
      registerTagMap_10_valid <= _GEN_857;
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_10_tagId <= 4'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      if (5'ha == io_decoders_0_destination_destinationRegister) begin // @[ReorderBuffer.scala 149:15]
        registerTagMap_10_tagId <= head; // @[ReorderBuffer.scala 149:15]
      end
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_11_valid <= 1'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      registerTagMap_11_valid <= _GEN_1405;
    end else if (canCommit_3) begin // @[ReorderBuffer.scala 88:21]
      if (_io_registerFile_3_valid_T) begin // @[ReorderBuffer.scala 89:22]
        registerTagMap_11_valid <= _GEN_1088;
      end else begin
        registerTagMap_11_valid <= _GEN_858;
      end
    end else begin
      registerTagMap_11_valid <= _GEN_858;
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_11_tagId <= 4'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      if (5'hb == io_decoders_0_destination_destinationRegister) begin // @[ReorderBuffer.scala 149:15]
        registerTagMap_11_tagId <= head; // @[ReorderBuffer.scala 149:15]
      end
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_12_valid <= 1'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      registerTagMap_12_valid <= _GEN_1406;
    end else if (canCommit_3) begin // @[ReorderBuffer.scala 88:21]
      if (_io_registerFile_3_valid_T) begin // @[ReorderBuffer.scala 89:22]
        registerTagMap_12_valid <= _GEN_1089;
      end else begin
        registerTagMap_12_valid <= _GEN_859;
      end
    end else begin
      registerTagMap_12_valid <= _GEN_859;
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_12_tagId <= 4'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      if (5'hc == io_decoders_0_destination_destinationRegister) begin // @[ReorderBuffer.scala 149:15]
        registerTagMap_12_tagId <= head; // @[ReorderBuffer.scala 149:15]
      end
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_13_valid <= 1'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      registerTagMap_13_valid <= _GEN_1407;
    end else if (canCommit_3) begin // @[ReorderBuffer.scala 88:21]
      if (_io_registerFile_3_valid_T) begin // @[ReorderBuffer.scala 89:22]
        registerTagMap_13_valid <= _GEN_1090;
      end else begin
        registerTagMap_13_valid <= _GEN_860;
      end
    end else begin
      registerTagMap_13_valid <= _GEN_860;
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_13_tagId <= 4'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      if (5'hd == io_decoders_0_destination_destinationRegister) begin // @[ReorderBuffer.scala 149:15]
        registerTagMap_13_tagId <= head; // @[ReorderBuffer.scala 149:15]
      end
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_14_valid <= 1'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      registerTagMap_14_valid <= _GEN_1408;
    end else if (canCommit_3) begin // @[ReorderBuffer.scala 88:21]
      if (_io_registerFile_3_valid_T) begin // @[ReorderBuffer.scala 89:22]
        registerTagMap_14_valid <= _GEN_1091;
      end else begin
        registerTagMap_14_valid <= _GEN_861;
      end
    end else begin
      registerTagMap_14_valid <= _GEN_861;
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_14_tagId <= 4'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      if (5'he == io_decoders_0_destination_destinationRegister) begin // @[ReorderBuffer.scala 149:15]
        registerTagMap_14_tagId <= head; // @[ReorderBuffer.scala 149:15]
      end
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_15_valid <= 1'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      registerTagMap_15_valid <= _GEN_1409;
    end else if (canCommit_3) begin // @[ReorderBuffer.scala 88:21]
      if (_io_registerFile_3_valid_T) begin // @[ReorderBuffer.scala 89:22]
        registerTagMap_15_valid <= _GEN_1092;
      end else begin
        registerTagMap_15_valid <= _GEN_862;
      end
    end else begin
      registerTagMap_15_valid <= _GEN_862;
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_15_tagId <= 4'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      if (5'hf == io_decoders_0_destination_destinationRegister) begin // @[ReorderBuffer.scala 149:15]
        registerTagMap_15_tagId <= head; // @[ReorderBuffer.scala 149:15]
      end
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_16_valid <= 1'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      registerTagMap_16_valid <= _GEN_1410;
    end else if (canCommit_3) begin // @[ReorderBuffer.scala 88:21]
      if (_io_registerFile_3_valid_T) begin // @[ReorderBuffer.scala 89:22]
        registerTagMap_16_valid <= _GEN_1093;
      end else begin
        registerTagMap_16_valid <= _GEN_863;
      end
    end else begin
      registerTagMap_16_valid <= _GEN_863;
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_16_tagId <= 4'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      if (5'h10 == io_decoders_0_destination_destinationRegister) begin // @[ReorderBuffer.scala 149:15]
        registerTagMap_16_tagId <= head; // @[ReorderBuffer.scala 149:15]
      end
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_17_valid <= 1'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      registerTagMap_17_valid <= _GEN_1411;
    end else if (canCommit_3) begin // @[ReorderBuffer.scala 88:21]
      if (_io_registerFile_3_valid_T) begin // @[ReorderBuffer.scala 89:22]
        registerTagMap_17_valid <= _GEN_1094;
      end else begin
        registerTagMap_17_valid <= _GEN_864;
      end
    end else begin
      registerTagMap_17_valid <= _GEN_864;
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_17_tagId <= 4'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      if (5'h11 == io_decoders_0_destination_destinationRegister) begin // @[ReorderBuffer.scala 149:15]
        registerTagMap_17_tagId <= head; // @[ReorderBuffer.scala 149:15]
      end
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_18_valid <= 1'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      registerTagMap_18_valid <= _GEN_1412;
    end else if (canCommit_3) begin // @[ReorderBuffer.scala 88:21]
      if (_io_registerFile_3_valid_T) begin // @[ReorderBuffer.scala 89:22]
        registerTagMap_18_valid <= _GEN_1095;
      end else begin
        registerTagMap_18_valid <= _GEN_865;
      end
    end else begin
      registerTagMap_18_valid <= _GEN_865;
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_18_tagId <= 4'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      if (5'h12 == io_decoders_0_destination_destinationRegister) begin // @[ReorderBuffer.scala 149:15]
        registerTagMap_18_tagId <= head; // @[ReorderBuffer.scala 149:15]
      end
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_19_valid <= 1'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      registerTagMap_19_valid <= _GEN_1413;
    end else if (canCommit_3) begin // @[ReorderBuffer.scala 88:21]
      if (_io_registerFile_3_valid_T) begin // @[ReorderBuffer.scala 89:22]
        registerTagMap_19_valid <= _GEN_1096;
      end else begin
        registerTagMap_19_valid <= _GEN_866;
      end
    end else begin
      registerTagMap_19_valid <= _GEN_866;
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_19_tagId <= 4'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      if (5'h13 == io_decoders_0_destination_destinationRegister) begin // @[ReorderBuffer.scala 149:15]
        registerTagMap_19_tagId <= head; // @[ReorderBuffer.scala 149:15]
      end
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_20_valid <= 1'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      registerTagMap_20_valid <= _GEN_1414;
    end else if (canCommit_3) begin // @[ReorderBuffer.scala 88:21]
      if (_io_registerFile_3_valid_T) begin // @[ReorderBuffer.scala 89:22]
        registerTagMap_20_valid <= _GEN_1097;
      end else begin
        registerTagMap_20_valid <= _GEN_867;
      end
    end else begin
      registerTagMap_20_valid <= _GEN_867;
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_20_tagId <= 4'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      if (5'h14 == io_decoders_0_destination_destinationRegister) begin // @[ReorderBuffer.scala 149:15]
        registerTagMap_20_tagId <= head; // @[ReorderBuffer.scala 149:15]
      end
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_21_valid <= 1'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      registerTagMap_21_valid <= _GEN_1415;
    end else if (canCommit_3) begin // @[ReorderBuffer.scala 88:21]
      if (_io_registerFile_3_valid_T) begin // @[ReorderBuffer.scala 89:22]
        registerTagMap_21_valid <= _GEN_1098;
      end else begin
        registerTagMap_21_valid <= _GEN_868;
      end
    end else begin
      registerTagMap_21_valid <= _GEN_868;
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_21_tagId <= 4'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      if (5'h15 == io_decoders_0_destination_destinationRegister) begin // @[ReorderBuffer.scala 149:15]
        registerTagMap_21_tagId <= head; // @[ReorderBuffer.scala 149:15]
      end
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_22_valid <= 1'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      registerTagMap_22_valid <= _GEN_1416;
    end else if (canCommit_3) begin // @[ReorderBuffer.scala 88:21]
      if (_io_registerFile_3_valid_T) begin // @[ReorderBuffer.scala 89:22]
        registerTagMap_22_valid <= _GEN_1099;
      end else begin
        registerTagMap_22_valid <= _GEN_869;
      end
    end else begin
      registerTagMap_22_valid <= _GEN_869;
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_22_tagId <= 4'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      if (5'h16 == io_decoders_0_destination_destinationRegister) begin // @[ReorderBuffer.scala 149:15]
        registerTagMap_22_tagId <= head; // @[ReorderBuffer.scala 149:15]
      end
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_23_valid <= 1'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      registerTagMap_23_valid <= _GEN_1417;
    end else if (canCommit_3) begin // @[ReorderBuffer.scala 88:21]
      if (_io_registerFile_3_valid_T) begin // @[ReorderBuffer.scala 89:22]
        registerTagMap_23_valid <= _GEN_1100;
      end else begin
        registerTagMap_23_valid <= _GEN_870;
      end
    end else begin
      registerTagMap_23_valid <= _GEN_870;
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_23_tagId <= 4'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      if (5'h17 == io_decoders_0_destination_destinationRegister) begin // @[ReorderBuffer.scala 149:15]
        registerTagMap_23_tagId <= head; // @[ReorderBuffer.scala 149:15]
      end
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_24_valid <= 1'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      registerTagMap_24_valid <= _GEN_1418;
    end else if (canCommit_3) begin // @[ReorderBuffer.scala 88:21]
      if (_io_registerFile_3_valid_T) begin // @[ReorderBuffer.scala 89:22]
        registerTagMap_24_valid <= _GEN_1101;
      end else begin
        registerTagMap_24_valid <= _GEN_871;
      end
    end else begin
      registerTagMap_24_valid <= _GEN_871;
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_24_tagId <= 4'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      if (5'h18 == io_decoders_0_destination_destinationRegister) begin // @[ReorderBuffer.scala 149:15]
        registerTagMap_24_tagId <= head; // @[ReorderBuffer.scala 149:15]
      end
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_25_valid <= 1'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      registerTagMap_25_valid <= _GEN_1419;
    end else if (canCommit_3) begin // @[ReorderBuffer.scala 88:21]
      if (_io_registerFile_3_valid_T) begin // @[ReorderBuffer.scala 89:22]
        registerTagMap_25_valid <= _GEN_1102;
      end else begin
        registerTagMap_25_valid <= _GEN_872;
      end
    end else begin
      registerTagMap_25_valid <= _GEN_872;
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_25_tagId <= 4'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      if (5'h19 == io_decoders_0_destination_destinationRegister) begin // @[ReorderBuffer.scala 149:15]
        registerTagMap_25_tagId <= head; // @[ReorderBuffer.scala 149:15]
      end
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_26_valid <= 1'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      registerTagMap_26_valid <= _GEN_1420;
    end else if (canCommit_3) begin // @[ReorderBuffer.scala 88:21]
      if (_io_registerFile_3_valid_T) begin // @[ReorderBuffer.scala 89:22]
        registerTagMap_26_valid <= _GEN_1103;
      end else begin
        registerTagMap_26_valid <= _GEN_873;
      end
    end else begin
      registerTagMap_26_valid <= _GEN_873;
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_26_tagId <= 4'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      if (5'h1a == io_decoders_0_destination_destinationRegister) begin // @[ReorderBuffer.scala 149:15]
        registerTagMap_26_tagId <= head; // @[ReorderBuffer.scala 149:15]
      end
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_27_valid <= 1'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      registerTagMap_27_valid <= _GEN_1421;
    end else if (canCommit_3) begin // @[ReorderBuffer.scala 88:21]
      if (_io_registerFile_3_valid_T) begin // @[ReorderBuffer.scala 89:22]
        registerTagMap_27_valid <= _GEN_1104;
      end else begin
        registerTagMap_27_valid <= _GEN_874;
      end
    end else begin
      registerTagMap_27_valid <= _GEN_874;
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_27_tagId <= 4'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      if (5'h1b == io_decoders_0_destination_destinationRegister) begin // @[ReorderBuffer.scala 149:15]
        registerTagMap_27_tagId <= head; // @[ReorderBuffer.scala 149:15]
      end
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_28_valid <= 1'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      registerTagMap_28_valid <= _GEN_1422;
    end else if (canCommit_3) begin // @[ReorderBuffer.scala 88:21]
      if (_io_registerFile_3_valid_T) begin // @[ReorderBuffer.scala 89:22]
        registerTagMap_28_valid <= _GEN_1105;
      end else begin
        registerTagMap_28_valid <= _GEN_875;
      end
    end else begin
      registerTagMap_28_valid <= _GEN_875;
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_28_tagId <= 4'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      if (5'h1c == io_decoders_0_destination_destinationRegister) begin // @[ReorderBuffer.scala 149:15]
        registerTagMap_28_tagId <= head; // @[ReorderBuffer.scala 149:15]
      end
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_29_valid <= 1'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      registerTagMap_29_valid <= _GEN_1423;
    end else if (canCommit_3) begin // @[ReorderBuffer.scala 88:21]
      if (_io_registerFile_3_valid_T) begin // @[ReorderBuffer.scala 89:22]
        registerTagMap_29_valid <= _GEN_1106;
      end else begin
        registerTagMap_29_valid <= _GEN_876;
      end
    end else begin
      registerTagMap_29_valid <= _GEN_876;
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_29_tagId <= 4'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      if (5'h1d == io_decoders_0_destination_destinationRegister) begin // @[ReorderBuffer.scala 149:15]
        registerTagMap_29_tagId <= head; // @[ReorderBuffer.scala 149:15]
      end
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_30_valid <= 1'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      registerTagMap_30_valid <= _GEN_1424;
    end else if (canCommit_3) begin // @[ReorderBuffer.scala 88:21]
      if (_io_registerFile_3_valid_T) begin // @[ReorderBuffer.scala 89:22]
        registerTagMap_30_valid <= _GEN_1107;
      end else begin
        registerTagMap_30_valid <= _GEN_877;
      end
    end else begin
      registerTagMap_30_valid <= _GEN_877;
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_30_tagId <= 4'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      if (5'h1e == io_decoders_0_destination_destinationRegister) begin // @[ReorderBuffer.scala 149:15]
        registerTagMap_30_tagId <= head; // @[ReorderBuffer.scala 149:15]
      end
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_31_valid <= 1'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      registerTagMap_31_valid <= _GEN_1425;
    end else if (canCommit_3) begin // @[ReorderBuffer.scala 88:21]
      if (_io_registerFile_3_valid_T) begin // @[ReorderBuffer.scala 89:22]
        registerTagMap_31_valid <= _GEN_1108;
      end else begin
        registerTagMap_31_valid <= _GEN_878;
      end
    end else begin
      registerTagMap_31_valid <= _GEN_878;
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_31_tagId <= 4'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      if (5'h1f == io_decoders_0_destination_destinationRegister) begin // @[ReorderBuffer.scala 149:15]
        registerTagMap_31_tagId <= head; // @[ReorderBuffer.scala 149:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  head = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  tail = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  buffer_0_destinationRegister = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  buffer_0_valueReady = _RAND_3[0:0];
  _RAND_4 = {2{`RANDOM}};
  buffer_0_value = _RAND_4[63:0];
  _RAND_5 = {1{`RANDOM}};
  buffer_0_storeSign = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  buffer_0_isError = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  buffer_1_destinationRegister = _RAND_7[4:0];
  _RAND_8 = {1{`RANDOM}};
  buffer_1_valueReady = _RAND_8[0:0];
  _RAND_9 = {2{`RANDOM}};
  buffer_1_value = _RAND_9[63:0];
  _RAND_10 = {1{`RANDOM}};
  buffer_1_storeSign = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  buffer_1_isError = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  buffer_2_destinationRegister = _RAND_12[4:0];
  _RAND_13 = {1{`RANDOM}};
  buffer_2_valueReady = _RAND_13[0:0];
  _RAND_14 = {2{`RANDOM}};
  buffer_2_value = _RAND_14[63:0];
  _RAND_15 = {1{`RANDOM}};
  buffer_2_storeSign = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  buffer_2_isError = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  buffer_3_destinationRegister = _RAND_17[4:0];
  _RAND_18 = {1{`RANDOM}};
  buffer_3_valueReady = _RAND_18[0:0];
  _RAND_19 = {2{`RANDOM}};
  buffer_3_value = _RAND_19[63:0];
  _RAND_20 = {1{`RANDOM}};
  buffer_3_storeSign = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  buffer_3_isError = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  buffer_4_destinationRegister = _RAND_22[4:0];
  _RAND_23 = {1{`RANDOM}};
  buffer_4_valueReady = _RAND_23[0:0];
  _RAND_24 = {2{`RANDOM}};
  buffer_4_value = _RAND_24[63:0];
  _RAND_25 = {1{`RANDOM}};
  buffer_4_storeSign = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  buffer_4_isError = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  buffer_5_destinationRegister = _RAND_27[4:0];
  _RAND_28 = {1{`RANDOM}};
  buffer_5_valueReady = _RAND_28[0:0];
  _RAND_29 = {2{`RANDOM}};
  buffer_5_value = _RAND_29[63:0];
  _RAND_30 = {1{`RANDOM}};
  buffer_5_storeSign = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  buffer_5_isError = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  buffer_6_destinationRegister = _RAND_32[4:0];
  _RAND_33 = {1{`RANDOM}};
  buffer_6_valueReady = _RAND_33[0:0];
  _RAND_34 = {2{`RANDOM}};
  buffer_6_value = _RAND_34[63:0];
  _RAND_35 = {1{`RANDOM}};
  buffer_6_storeSign = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  buffer_6_isError = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  buffer_7_destinationRegister = _RAND_37[4:0];
  _RAND_38 = {1{`RANDOM}};
  buffer_7_valueReady = _RAND_38[0:0];
  _RAND_39 = {2{`RANDOM}};
  buffer_7_value = _RAND_39[63:0];
  _RAND_40 = {1{`RANDOM}};
  buffer_7_storeSign = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  buffer_7_isError = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  buffer_8_destinationRegister = _RAND_42[4:0];
  _RAND_43 = {1{`RANDOM}};
  buffer_8_valueReady = _RAND_43[0:0];
  _RAND_44 = {2{`RANDOM}};
  buffer_8_value = _RAND_44[63:0];
  _RAND_45 = {1{`RANDOM}};
  buffer_8_storeSign = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  buffer_8_isError = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  buffer_9_destinationRegister = _RAND_47[4:0];
  _RAND_48 = {1{`RANDOM}};
  buffer_9_valueReady = _RAND_48[0:0];
  _RAND_49 = {2{`RANDOM}};
  buffer_9_value = _RAND_49[63:0];
  _RAND_50 = {1{`RANDOM}};
  buffer_9_storeSign = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  buffer_9_isError = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  buffer_10_destinationRegister = _RAND_52[4:0];
  _RAND_53 = {1{`RANDOM}};
  buffer_10_valueReady = _RAND_53[0:0];
  _RAND_54 = {2{`RANDOM}};
  buffer_10_value = _RAND_54[63:0];
  _RAND_55 = {1{`RANDOM}};
  buffer_10_storeSign = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  buffer_10_isError = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  buffer_11_destinationRegister = _RAND_57[4:0];
  _RAND_58 = {1{`RANDOM}};
  buffer_11_valueReady = _RAND_58[0:0];
  _RAND_59 = {2{`RANDOM}};
  buffer_11_value = _RAND_59[63:0];
  _RAND_60 = {1{`RANDOM}};
  buffer_11_storeSign = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  buffer_11_isError = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  buffer_12_destinationRegister = _RAND_62[4:0];
  _RAND_63 = {1{`RANDOM}};
  buffer_12_valueReady = _RAND_63[0:0];
  _RAND_64 = {2{`RANDOM}};
  buffer_12_value = _RAND_64[63:0];
  _RAND_65 = {1{`RANDOM}};
  buffer_12_storeSign = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  buffer_12_isError = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  buffer_13_destinationRegister = _RAND_67[4:0];
  _RAND_68 = {1{`RANDOM}};
  buffer_13_valueReady = _RAND_68[0:0];
  _RAND_69 = {2{`RANDOM}};
  buffer_13_value = _RAND_69[63:0];
  _RAND_70 = {1{`RANDOM}};
  buffer_13_storeSign = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  buffer_13_isError = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  buffer_14_destinationRegister = _RAND_72[4:0];
  _RAND_73 = {1{`RANDOM}};
  buffer_14_valueReady = _RAND_73[0:0];
  _RAND_74 = {2{`RANDOM}};
  buffer_14_value = _RAND_74[63:0];
  _RAND_75 = {1{`RANDOM}};
  buffer_14_storeSign = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  buffer_14_isError = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  buffer_15_destinationRegister = _RAND_77[4:0];
  _RAND_78 = {1{`RANDOM}};
  buffer_15_valueReady = _RAND_78[0:0];
  _RAND_79 = {2{`RANDOM}};
  buffer_15_value = _RAND_79[63:0];
  _RAND_80 = {1{`RANDOM}};
  buffer_15_storeSign = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  buffer_15_isError = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  registerTagMap_1_valid = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  registerTagMap_1_tagId = _RAND_83[3:0];
  _RAND_84 = {1{`RANDOM}};
  registerTagMap_2_valid = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  registerTagMap_2_tagId = _RAND_85[3:0];
  _RAND_86 = {1{`RANDOM}};
  registerTagMap_3_valid = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  registerTagMap_3_tagId = _RAND_87[3:0];
  _RAND_88 = {1{`RANDOM}};
  registerTagMap_4_valid = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  registerTagMap_4_tagId = _RAND_89[3:0];
  _RAND_90 = {1{`RANDOM}};
  registerTagMap_5_valid = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  registerTagMap_5_tagId = _RAND_91[3:0];
  _RAND_92 = {1{`RANDOM}};
  registerTagMap_6_valid = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  registerTagMap_6_tagId = _RAND_93[3:0];
  _RAND_94 = {1{`RANDOM}};
  registerTagMap_7_valid = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  registerTagMap_7_tagId = _RAND_95[3:0];
  _RAND_96 = {1{`RANDOM}};
  registerTagMap_8_valid = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  registerTagMap_8_tagId = _RAND_97[3:0];
  _RAND_98 = {1{`RANDOM}};
  registerTagMap_9_valid = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  registerTagMap_9_tagId = _RAND_99[3:0];
  _RAND_100 = {1{`RANDOM}};
  registerTagMap_10_valid = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  registerTagMap_10_tagId = _RAND_101[3:0];
  _RAND_102 = {1{`RANDOM}};
  registerTagMap_11_valid = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  registerTagMap_11_tagId = _RAND_103[3:0];
  _RAND_104 = {1{`RANDOM}};
  registerTagMap_12_valid = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  registerTagMap_12_tagId = _RAND_105[3:0];
  _RAND_106 = {1{`RANDOM}};
  registerTagMap_13_valid = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  registerTagMap_13_tagId = _RAND_107[3:0];
  _RAND_108 = {1{`RANDOM}};
  registerTagMap_14_valid = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  registerTagMap_14_tagId = _RAND_109[3:0];
  _RAND_110 = {1{`RANDOM}};
  registerTagMap_15_valid = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  registerTagMap_15_tagId = _RAND_111[3:0];
  _RAND_112 = {1{`RANDOM}};
  registerTagMap_16_valid = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  registerTagMap_16_tagId = _RAND_113[3:0];
  _RAND_114 = {1{`RANDOM}};
  registerTagMap_17_valid = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  registerTagMap_17_tagId = _RAND_115[3:0];
  _RAND_116 = {1{`RANDOM}};
  registerTagMap_18_valid = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  registerTagMap_18_tagId = _RAND_117[3:0];
  _RAND_118 = {1{`RANDOM}};
  registerTagMap_19_valid = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  registerTagMap_19_tagId = _RAND_119[3:0];
  _RAND_120 = {1{`RANDOM}};
  registerTagMap_20_valid = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  registerTagMap_20_tagId = _RAND_121[3:0];
  _RAND_122 = {1{`RANDOM}};
  registerTagMap_21_valid = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  registerTagMap_21_tagId = _RAND_123[3:0];
  _RAND_124 = {1{`RANDOM}};
  registerTagMap_22_valid = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  registerTagMap_22_tagId = _RAND_125[3:0];
  _RAND_126 = {1{`RANDOM}};
  registerTagMap_23_valid = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  registerTagMap_23_tagId = _RAND_127[3:0];
  _RAND_128 = {1{`RANDOM}};
  registerTagMap_24_valid = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  registerTagMap_24_tagId = _RAND_129[3:0];
  _RAND_130 = {1{`RANDOM}};
  registerTagMap_25_valid = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  registerTagMap_25_tagId = _RAND_131[3:0];
  _RAND_132 = {1{`RANDOM}};
  registerTagMap_26_valid = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  registerTagMap_26_tagId = _RAND_133[3:0];
  _RAND_134 = {1{`RANDOM}};
  registerTagMap_27_valid = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  registerTagMap_27_tagId = _RAND_135[3:0];
  _RAND_136 = {1{`RANDOM}};
  registerTagMap_28_valid = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  registerTagMap_28_tagId = _RAND_137[3:0];
  _RAND_138 = {1{`RANDOM}};
  registerTagMap_29_valid = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  registerTagMap_29_tagId = _RAND_139[3:0];
  _RAND_140 = {1{`RANDOM}};
  registerTagMap_30_valid = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  registerTagMap_30_tagId = _RAND_141[3:0];
  _RAND_142 = {1{`RANDOM}};
  registerTagMap_31_valid = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  registerTagMap_31_tagId = _RAND_143[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ReorderBuffer_1(
  input         clock,
  input         reset,
  input  [4:0]  io_decoders_0_source1_sourceRegister,
  output        io_decoders_0_source1_matchingTag_valid,
  output [3:0]  io_decoders_0_source1_matchingTag_bits_id,
  output        io_decoders_0_source1_value_valid,
  output [63:0] io_decoders_0_source1_value_bits,
  input  [4:0]  io_decoders_0_source2_sourceRegister,
  output        io_decoders_0_source2_matchingTag_valid,
  output [3:0]  io_decoders_0_source2_matchingTag_bits_id,
  output        io_decoders_0_source2_value_valid,
  output [63:0] io_decoders_0_source2_value_bits,
  input  [4:0]  io_decoders_0_destination_destinationRegister,
  output [3:0]  io_decoders_0_destination_destinationTag_id,
  input         io_decoders_0_destination_storeSign,
  output        io_decoders_0_ready,
  input         io_decoders_0_valid,
  input         io_collectedOutputs_outputs_valid,
  input         io_collectedOutputs_outputs_bits_resultType,
  input  [63:0] io_collectedOutputs_outputs_bits_value,
  input         io_collectedOutputs_outputs_bits_isError,
  input         io_collectedOutputs_outputs_bits_tag_threadId,
  input  [3:0]  io_collectedOutputs_outputs_bits_tag_id,
  output        io_registerFile_0_valid,
  output [4:0]  io_registerFile_0_bits_destinationRegister,
  output [63:0] io_registerFile_0_bits_value,
  output        io_registerFile_1_valid,
  output [4:0]  io_registerFile_1_bits_destinationRegister,
  output [63:0] io_registerFile_1_bits_value,
  output        io_registerFile_2_valid,
  output [4:0]  io_registerFile_2_bits_destinationRegister,
  output [63:0] io_registerFile_2_bits_value,
  output        io_registerFile_3_valid,
  output [4:0]  io_registerFile_3_bits_destinationRegister,
  output [63:0] io_registerFile_3_bits_value,
  output        io_loadStoreQueue_0_valid,
  output [3:0]  io_loadStoreQueue_0_bits_destinationTag_id,
  output        io_loadStoreQueue_1_valid,
  output [3:0]  io_loadStoreQueue_1_bits_destinationTag_id,
  output        io_loadStoreQueue_2_valid,
  output [3:0]  io_loadStoreQueue_2_bits_destinationTag_id,
  output        io_loadStoreQueue_3_valid,
  output [3:0]  io_loadStoreQueue_3_bits_destinationTag_id,
  output        io_isEmpty,
  output [1:0]  io_csr_retireCount,
  output        io_isError
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [63:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [63:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [63:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [63:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [63:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [63:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [63:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [63:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] head; // @[ReorderBuffer.scala 53:21]
  reg [3:0] tail; // @[ReorderBuffer.scala 54:21]
  reg [4:0] buffer_0_destinationRegister; // @[ReorderBuffer.scala 55:23]
  reg  buffer_0_valueReady; // @[ReorderBuffer.scala 55:23]
  reg [63:0] buffer_0_value; // @[ReorderBuffer.scala 55:23]
  reg  buffer_0_storeSign; // @[ReorderBuffer.scala 55:23]
  reg  buffer_0_isError; // @[ReorderBuffer.scala 55:23]
  reg [4:0] buffer_1_destinationRegister; // @[ReorderBuffer.scala 55:23]
  reg  buffer_1_valueReady; // @[ReorderBuffer.scala 55:23]
  reg [63:0] buffer_1_value; // @[ReorderBuffer.scala 55:23]
  reg  buffer_1_storeSign; // @[ReorderBuffer.scala 55:23]
  reg  buffer_1_isError; // @[ReorderBuffer.scala 55:23]
  reg [4:0] buffer_2_destinationRegister; // @[ReorderBuffer.scala 55:23]
  reg  buffer_2_valueReady; // @[ReorderBuffer.scala 55:23]
  reg [63:0] buffer_2_value; // @[ReorderBuffer.scala 55:23]
  reg  buffer_2_storeSign; // @[ReorderBuffer.scala 55:23]
  reg  buffer_2_isError; // @[ReorderBuffer.scala 55:23]
  reg [4:0] buffer_3_destinationRegister; // @[ReorderBuffer.scala 55:23]
  reg  buffer_3_valueReady; // @[ReorderBuffer.scala 55:23]
  reg [63:0] buffer_3_value; // @[ReorderBuffer.scala 55:23]
  reg  buffer_3_storeSign; // @[ReorderBuffer.scala 55:23]
  reg  buffer_3_isError; // @[ReorderBuffer.scala 55:23]
  reg [4:0] buffer_4_destinationRegister; // @[ReorderBuffer.scala 55:23]
  reg  buffer_4_valueReady; // @[ReorderBuffer.scala 55:23]
  reg [63:0] buffer_4_value; // @[ReorderBuffer.scala 55:23]
  reg  buffer_4_storeSign; // @[ReorderBuffer.scala 55:23]
  reg  buffer_4_isError; // @[ReorderBuffer.scala 55:23]
  reg [4:0] buffer_5_destinationRegister; // @[ReorderBuffer.scala 55:23]
  reg  buffer_5_valueReady; // @[ReorderBuffer.scala 55:23]
  reg [63:0] buffer_5_value; // @[ReorderBuffer.scala 55:23]
  reg  buffer_5_storeSign; // @[ReorderBuffer.scala 55:23]
  reg  buffer_5_isError; // @[ReorderBuffer.scala 55:23]
  reg [4:0] buffer_6_destinationRegister; // @[ReorderBuffer.scala 55:23]
  reg  buffer_6_valueReady; // @[ReorderBuffer.scala 55:23]
  reg [63:0] buffer_6_value; // @[ReorderBuffer.scala 55:23]
  reg  buffer_6_storeSign; // @[ReorderBuffer.scala 55:23]
  reg  buffer_6_isError; // @[ReorderBuffer.scala 55:23]
  reg [4:0] buffer_7_destinationRegister; // @[ReorderBuffer.scala 55:23]
  reg  buffer_7_valueReady; // @[ReorderBuffer.scala 55:23]
  reg [63:0] buffer_7_value; // @[ReorderBuffer.scala 55:23]
  reg  buffer_7_storeSign; // @[ReorderBuffer.scala 55:23]
  reg  buffer_7_isError; // @[ReorderBuffer.scala 55:23]
  reg [4:0] buffer_8_destinationRegister; // @[ReorderBuffer.scala 55:23]
  reg  buffer_8_valueReady; // @[ReorderBuffer.scala 55:23]
  reg [63:0] buffer_8_value; // @[ReorderBuffer.scala 55:23]
  reg  buffer_8_storeSign; // @[ReorderBuffer.scala 55:23]
  reg  buffer_8_isError; // @[ReorderBuffer.scala 55:23]
  reg [4:0] buffer_9_destinationRegister; // @[ReorderBuffer.scala 55:23]
  reg  buffer_9_valueReady; // @[ReorderBuffer.scala 55:23]
  reg [63:0] buffer_9_value; // @[ReorderBuffer.scala 55:23]
  reg  buffer_9_storeSign; // @[ReorderBuffer.scala 55:23]
  reg  buffer_9_isError; // @[ReorderBuffer.scala 55:23]
  reg [4:0] buffer_10_destinationRegister; // @[ReorderBuffer.scala 55:23]
  reg  buffer_10_valueReady; // @[ReorderBuffer.scala 55:23]
  reg [63:0] buffer_10_value; // @[ReorderBuffer.scala 55:23]
  reg  buffer_10_storeSign; // @[ReorderBuffer.scala 55:23]
  reg  buffer_10_isError; // @[ReorderBuffer.scala 55:23]
  reg [4:0] buffer_11_destinationRegister; // @[ReorderBuffer.scala 55:23]
  reg  buffer_11_valueReady; // @[ReorderBuffer.scala 55:23]
  reg [63:0] buffer_11_value; // @[ReorderBuffer.scala 55:23]
  reg  buffer_11_storeSign; // @[ReorderBuffer.scala 55:23]
  reg  buffer_11_isError; // @[ReorderBuffer.scala 55:23]
  reg [4:0] buffer_12_destinationRegister; // @[ReorderBuffer.scala 55:23]
  reg  buffer_12_valueReady; // @[ReorderBuffer.scala 55:23]
  reg [63:0] buffer_12_value; // @[ReorderBuffer.scala 55:23]
  reg  buffer_12_storeSign; // @[ReorderBuffer.scala 55:23]
  reg  buffer_12_isError; // @[ReorderBuffer.scala 55:23]
  reg [4:0] buffer_13_destinationRegister; // @[ReorderBuffer.scala 55:23]
  reg  buffer_13_valueReady; // @[ReorderBuffer.scala 55:23]
  reg [63:0] buffer_13_value; // @[ReorderBuffer.scala 55:23]
  reg  buffer_13_storeSign; // @[ReorderBuffer.scala 55:23]
  reg  buffer_13_isError; // @[ReorderBuffer.scala 55:23]
  reg [4:0] buffer_14_destinationRegister; // @[ReorderBuffer.scala 55:23]
  reg  buffer_14_valueReady; // @[ReorderBuffer.scala 55:23]
  reg [63:0] buffer_14_value; // @[ReorderBuffer.scala 55:23]
  reg  buffer_14_storeSign; // @[ReorderBuffer.scala 55:23]
  reg  buffer_14_isError; // @[ReorderBuffer.scala 55:23]
  reg [4:0] buffer_15_destinationRegister; // @[ReorderBuffer.scala 55:23]
  reg  buffer_15_valueReady; // @[ReorderBuffer.scala 55:23]
  reg [63:0] buffer_15_value; // @[ReorderBuffer.scala 55:23]
  reg  buffer_15_storeSign; // @[ReorderBuffer.scala 55:23]
  reg  buffer_15_isError; // @[ReorderBuffer.scala 55:23]
  reg  registerTagMap_1_valid; // @[ReorderBuffer.scala 69:39]
  reg [3:0] registerTagMap_1_tagId; // @[ReorderBuffer.scala 69:39]
  reg  registerTagMap_2_valid; // @[ReorderBuffer.scala 69:39]
  reg [3:0] registerTagMap_2_tagId; // @[ReorderBuffer.scala 69:39]
  reg  registerTagMap_3_valid; // @[ReorderBuffer.scala 69:39]
  reg [3:0] registerTagMap_3_tagId; // @[ReorderBuffer.scala 69:39]
  reg  registerTagMap_4_valid; // @[ReorderBuffer.scala 69:39]
  reg [3:0] registerTagMap_4_tagId; // @[ReorderBuffer.scala 69:39]
  reg  registerTagMap_5_valid; // @[ReorderBuffer.scala 69:39]
  reg [3:0] registerTagMap_5_tagId; // @[ReorderBuffer.scala 69:39]
  reg  registerTagMap_6_valid; // @[ReorderBuffer.scala 69:39]
  reg [3:0] registerTagMap_6_tagId; // @[ReorderBuffer.scala 69:39]
  reg  registerTagMap_7_valid; // @[ReorderBuffer.scala 69:39]
  reg [3:0] registerTagMap_7_tagId; // @[ReorderBuffer.scala 69:39]
  reg  registerTagMap_8_valid; // @[ReorderBuffer.scala 69:39]
  reg [3:0] registerTagMap_8_tagId; // @[ReorderBuffer.scala 69:39]
  reg  registerTagMap_9_valid; // @[ReorderBuffer.scala 69:39]
  reg [3:0] registerTagMap_9_tagId; // @[ReorderBuffer.scala 69:39]
  reg  registerTagMap_10_valid; // @[ReorderBuffer.scala 69:39]
  reg [3:0] registerTagMap_10_tagId; // @[ReorderBuffer.scala 69:39]
  reg  registerTagMap_11_valid; // @[ReorderBuffer.scala 69:39]
  reg [3:0] registerTagMap_11_tagId; // @[ReorderBuffer.scala 69:39]
  reg  registerTagMap_12_valid; // @[ReorderBuffer.scala 69:39]
  reg [3:0] registerTagMap_12_tagId; // @[ReorderBuffer.scala 69:39]
  reg  registerTagMap_13_valid; // @[ReorderBuffer.scala 69:39]
  reg [3:0] registerTagMap_13_tagId; // @[ReorderBuffer.scala 69:39]
  reg  registerTagMap_14_valid; // @[ReorderBuffer.scala 69:39]
  reg [3:0] registerTagMap_14_tagId; // @[ReorderBuffer.scala 69:39]
  reg  registerTagMap_15_valid; // @[ReorderBuffer.scala 69:39]
  reg [3:0] registerTagMap_15_tagId; // @[ReorderBuffer.scala 69:39]
  reg  registerTagMap_16_valid; // @[ReorderBuffer.scala 69:39]
  reg [3:0] registerTagMap_16_tagId; // @[ReorderBuffer.scala 69:39]
  reg  registerTagMap_17_valid; // @[ReorderBuffer.scala 69:39]
  reg [3:0] registerTagMap_17_tagId; // @[ReorderBuffer.scala 69:39]
  reg  registerTagMap_18_valid; // @[ReorderBuffer.scala 69:39]
  reg [3:0] registerTagMap_18_tagId; // @[ReorderBuffer.scala 69:39]
  reg  registerTagMap_19_valid; // @[ReorderBuffer.scala 69:39]
  reg [3:0] registerTagMap_19_tagId; // @[ReorderBuffer.scala 69:39]
  reg  registerTagMap_20_valid; // @[ReorderBuffer.scala 69:39]
  reg [3:0] registerTagMap_20_tagId; // @[ReorderBuffer.scala 69:39]
  reg  registerTagMap_21_valid; // @[ReorderBuffer.scala 69:39]
  reg [3:0] registerTagMap_21_tagId; // @[ReorderBuffer.scala 69:39]
  reg  registerTagMap_22_valid; // @[ReorderBuffer.scala 69:39]
  reg [3:0] registerTagMap_22_tagId; // @[ReorderBuffer.scala 69:39]
  reg  registerTagMap_23_valid; // @[ReorderBuffer.scala 69:39]
  reg [3:0] registerTagMap_23_tagId; // @[ReorderBuffer.scala 69:39]
  reg  registerTagMap_24_valid; // @[ReorderBuffer.scala 69:39]
  reg [3:0] registerTagMap_24_tagId; // @[ReorderBuffer.scala 69:39]
  reg  registerTagMap_25_valid; // @[ReorderBuffer.scala 69:39]
  reg [3:0] registerTagMap_25_tagId; // @[ReorderBuffer.scala 69:39]
  reg  registerTagMap_26_valid; // @[ReorderBuffer.scala 69:39]
  reg [3:0] registerTagMap_26_tagId; // @[ReorderBuffer.scala 69:39]
  reg  registerTagMap_27_valid; // @[ReorderBuffer.scala 69:39]
  reg [3:0] registerTagMap_27_tagId; // @[ReorderBuffer.scala 69:39]
  reg  registerTagMap_28_valid; // @[ReorderBuffer.scala 69:39]
  reg [3:0] registerTagMap_28_tagId; // @[ReorderBuffer.scala 69:39]
  reg  registerTagMap_29_valid; // @[ReorderBuffer.scala 69:39]
  reg [3:0] registerTagMap_29_tagId; // @[ReorderBuffer.scala 69:39]
  reg  registerTagMap_30_valid; // @[ReorderBuffer.scala 69:39]
  reg [3:0] registerTagMap_30_tagId; // @[ReorderBuffer.scala 69:39]
  reg  registerTagMap_31_valid; // @[ReorderBuffer.scala 69:39]
  reg [3:0] registerTagMap_31_tagId; // @[ReorderBuffer.scala 69:39]
  wire [4:0] _index_T = {{1'd0}, tail}; // @[ReorderBuffer.scala 77:22]
  wire [3:0] index = _index_T[3:0]; // @[ReorderBuffer.scala 77:22]
  wire  _GEN_1 = 4'h1 == index ? buffer_1_valueReady : buffer_0_valueReady; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_2 = 4'h2 == index ? buffer_2_valueReady : _GEN_1; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_3 = 4'h3 == index ? buffer_3_valueReady : _GEN_2; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_4 = 4'h4 == index ? buffer_4_valueReady : _GEN_3; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_5 = 4'h5 == index ? buffer_5_valueReady : _GEN_4; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_6 = 4'h6 == index ? buffer_6_valueReady : _GEN_5; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_7 = 4'h7 == index ? buffer_7_valueReady : _GEN_6; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_8 = 4'h8 == index ? buffer_8_valueReady : _GEN_7; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_9 = 4'h9 == index ? buffer_9_valueReady : _GEN_8; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_10 = 4'ha == index ? buffer_10_valueReady : _GEN_9; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_11 = 4'hb == index ? buffer_11_valueReady : _GEN_10; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_12 = 4'hc == index ? buffer_12_valueReady : _GEN_11; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_13 = 4'hd == index ? buffer_13_valueReady : _GEN_12; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_14 = 4'he == index ? buffer_14_valueReady : _GEN_13; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_15 = 4'hf == index ? buffer_15_valueReady : _GEN_14; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_17 = 4'h1 == index ? buffer_1_storeSign : buffer_0_storeSign; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_18 = 4'h2 == index ? buffer_2_storeSign : _GEN_17; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_19 = 4'h3 == index ? buffer_3_storeSign : _GEN_18; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_20 = 4'h4 == index ? buffer_4_storeSign : _GEN_19; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_21 = 4'h5 == index ? buffer_5_storeSign : _GEN_20; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_22 = 4'h6 == index ? buffer_6_storeSign : _GEN_21; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_23 = 4'h7 == index ? buffer_7_storeSign : _GEN_22; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_24 = 4'h8 == index ? buffer_8_storeSign : _GEN_23; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_25 = 4'h9 == index ? buffer_9_storeSign : _GEN_24; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_26 = 4'ha == index ? buffer_10_storeSign : _GEN_25; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_27 = 4'hb == index ? buffer_11_storeSign : _GEN_26; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_28 = 4'hc == index ? buffer_12_storeSign : _GEN_27; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_29 = 4'hd == index ? buffer_13_storeSign : _GEN_28; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_30 = 4'he == index ? buffer_14_storeSign : _GEN_29; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_31 = 4'hf == index ? buffer_15_storeSign : _GEN_30; // @[ReorderBuffer.scala 79:{50,50}]
  wire  instructionOk = _GEN_15 | _GEN_31; // @[ReorderBuffer.scala 79:50]
  wire  canCommit = index != head & instructionOk; // @[ReorderBuffer.scala 80:49]
  wire  _GEN_33 = 4'h1 == index ? buffer_1_isError : buffer_0_isError; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_34 = 4'h2 == index ? buffer_2_isError : _GEN_33; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_35 = 4'h3 == index ? buffer_3_isError : _GEN_34; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_36 = 4'h4 == index ? buffer_4_isError : _GEN_35; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_37 = 4'h5 == index ? buffer_5_isError : _GEN_36; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_38 = 4'h6 == index ? buffer_6_isError : _GEN_37; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_39 = 4'h7 == index ? buffer_7_isError : _GEN_38; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_40 = 4'h8 == index ? buffer_8_isError : _GEN_39; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_41 = 4'h9 == index ? buffer_9_isError : _GEN_40; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_42 = 4'ha == index ? buffer_10_isError : _GEN_41; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_43 = 4'hb == index ? buffer_11_isError : _GEN_42; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_44 = 4'hc == index ? buffer_12_isError : _GEN_43; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_45 = 4'hd == index ? buffer_13_isError : _GEN_44; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_46 = 4'he == index ? buffer_14_isError : _GEN_45; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_47 = 4'hf == index ? buffer_15_isError : _GEN_46; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _io_registerFile_0_valid_T = ~_GEN_47; // @[ReorderBuffer.scala 83:30]
  wire [63:0] _GEN_49 = 4'h1 == index ? buffer_1_value : buffer_0_value; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_50 = 4'h2 == index ? buffer_2_value : _GEN_49; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_51 = 4'h3 == index ? buffer_3_value : _GEN_50; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_52 = 4'h4 == index ? buffer_4_value : _GEN_51; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_53 = 4'h5 == index ? buffer_5_value : _GEN_52; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_54 = 4'h6 == index ? buffer_6_value : _GEN_53; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_55 = 4'h7 == index ? buffer_7_value : _GEN_54; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_56 = 4'h8 == index ? buffer_8_value : _GEN_55; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_57 = 4'h9 == index ? buffer_9_value : _GEN_56; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_58 = 4'ha == index ? buffer_10_value : _GEN_57; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_59 = 4'hb == index ? buffer_11_value : _GEN_58; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_60 = 4'hc == index ? buffer_12_value : _GEN_59; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_61 = 4'hd == index ? buffer_13_value : _GEN_60; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_62 = 4'he == index ? buffer_14_value : _GEN_61; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_63 = 4'hf == index ? buffer_15_value : _GEN_62; // @[ReorderBuffer.scala 90:{23,23}]
  wire [4:0] _GEN_65 = 4'h1 == index ? buffer_1_destinationRegister : buffer_0_destinationRegister; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_66 = 4'h2 == index ? buffer_2_destinationRegister : _GEN_65; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_67 = 4'h3 == index ? buffer_3_destinationRegister : _GEN_66; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_68 = 4'h4 == index ? buffer_4_destinationRegister : _GEN_67; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_69 = 4'h5 == index ? buffer_5_destinationRegister : _GEN_68; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_70 = 4'h6 == index ? buffer_6_destinationRegister : _GEN_69; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_71 = 4'h7 == index ? buffer_7_destinationRegister : _GEN_70; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_72 = 4'h8 == index ? buffer_8_destinationRegister : _GEN_71; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_73 = 4'h9 == index ? buffer_9_destinationRegister : _GEN_72; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_74 = 4'ha == index ? buffer_10_destinationRegister : _GEN_73; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_75 = 4'hb == index ? buffer_11_destinationRegister : _GEN_74; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_76 = 4'hc == index ? buffer_12_destinationRegister : _GEN_75; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_77 = 4'hd == index ? buffer_13_destinationRegister : _GEN_76; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_78 = 4'he == index ? buffer_14_destinationRegister : _GEN_77; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_79 = 4'hf == index ? buffer_15_destinationRegister : _GEN_78; // @[ReorderBuffer.scala 91:{37,37}]
  wire [3:0] _GEN_81 = 5'h1 == _GEN_79 ? registerTagMap_1_tagId : 4'h0; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_82 = 5'h2 == _GEN_79 ? registerTagMap_2_tagId : _GEN_81; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_83 = 5'h3 == _GEN_79 ? registerTagMap_3_tagId : _GEN_82; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_84 = 5'h4 == _GEN_79 ? registerTagMap_4_tagId : _GEN_83; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_85 = 5'h5 == _GEN_79 ? registerTagMap_5_tagId : _GEN_84; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_86 = 5'h6 == _GEN_79 ? registerTagMap_6_tagId : _GEN_85; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_87 = 5'h7 == _GEN_79 ? registerTagMap_7_tagId : _GEN_86; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_88 = 5'h8 == _GEN_79 ? registerTagMap_8_tagId : _GEN_87; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_89 = 5'h9 == _GEN_79 ? registerTagMap_9_tagId : _GEN_88; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_90 = 5'ha == _GEN_79 ? registerTagMap_10_tagId : _GEN_89; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_91 = 5'hb == _GEN_79 ? registerTagMap_11_tagId : _GEN_90; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_92 = 5'hc == _GEN_79 ? registerTagMap_12_tagId : _GEN_91; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_93 = 5'hd == _GEN_79 ? registerTagMap_13_tagId : _GEN_92; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_94 = 5'he == _GEN_79 ? registerTagMap_14_tagId : _GEN_93; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_95 = 5'hf == _GEN_79 ? registerTagMap_15_tagId : _GEN_94; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_96 = 5'h10 == _GEN_79 ? registerTagMap_16_tagId : _GEN_95; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_97 = 5'h11 == _GEN_79 ? registerTagMap_17_tagId : _GEN_96; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_98 = 5'h12 == _GEN_79 ? registerTagMap_18_tagId : _GEN_97; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_99 = 5'h13 == _GEN_79 ? registerTagMap_19_tagId : _GEN_98; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_100 = 5'h14 == _GEN_79 ? registerTagMap_20_tagId : _GEN_99; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_101 = 5'h15 == _GEN_79 ? registerTagMap_21_tagId : _GEN_100; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_102 = 5'h16 == _GEN_79 ? registerTagMap_22_tagId : _GEN_101; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_103 = 5'h17 == _GEN_79 ? registerTagMap_23_tagId : _GEN_102; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_104 = 5'h18 == _GEN_79 ? registerTagMap_24_tagId : _GEN_103; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_105 = 5'h19 == _GEN_79 ? registerTagMap_25_tagId : _GEN_104; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_106 = 5'h1a == _GEN_79 ? registerTagMap_26_tagId : _GEN_105; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_107 = 5'h1b == _GEN_79 ? registerTagMap_27_tagId : _GEN_106; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_108 = 5'h1c == _GEN_79 ? registerTagMap_28_tagId : _GEN_107; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_109 = 5'h1d == _GEN_79 ? registerTagMap_29_tagId : _GEN_108; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_110 = 5'h1e == _GEN_79 ? registerTagMap_30_tagId : _GEN_109; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_111 = 5'h1f == _GEN_79 ? registerTagMap_31_tagId : _GEN_110; // @[ReorderBuffer.scala 93:{17,17}]
  wire  _T_1 = index == _GEN_111; // @[ReorderBuffer.scala 93:17]
  wire  _GEN_145 = 5'h1 == _GEN_79 ? 1'h0 : registerTagMap_1_valid; // @[ReorderBuffer.scala 97:{13,13} 69:39]
  wire  _GEN_146 = 5'h2 == _GEN_79 ? 1'h0 : registerTagMap_2_valid; // @[ReorderBuffer.scala 97:{13,13} 69:39]
  wire  _GEN_147 = 5'h3 == _GEN_79 ? 1'h0 : registerTagMap_3_valid; // @[ReorderBuffer.scala 97:{13,13} 69:39]
  wire  _GEN_148 = 5'h4 == _GEN_79 ? 1'h0 : registerTagMap_4_valid; // @[ReorderBuffer.scala 97:{13,13} 69:39]
  wire  _GEN_149 = 5'h5 == _GEN_79 ? 1'h0 : registerTagMap_5_valid; // @[ReorderBuffer.scala 97:{13,13} 69:39]
  wire  _GEN_150 = 5'h6 == _GEN_79 ? 1'h0 : registerTagMap_6_valid; // @[ReorderBuffer.scala 97:{13,13} 69:39]
  wire  _GEN_151 = 5'h7 == _GEN_79 ? 1'h0 : registerTagMap_7_valid; // @[ReorderBuffer.scala 97:{13,13} 69:39]
  wire  _GEN_152 = 5'h8 == _GEN_79 ? 1'h0 : registerTagMap_8_valid; // @[ReorderBuffer.scala 97:{13,13} 69:39]
  wire  _GEN_153 = 5'h9 == _GEN_79 ? 1'h0 : registerTagMap_9_valid; // @[ReorderBuffer.scala 97:{13,13} 69:39]
  wire  _GEN_154 = 5'ha == _GEN_79 ? 1'h0 : registerTagMap_10_valid; // @[ReorderBuffer.scala 97:{13,13} 69:39]
  wire  _GEN_155 = 5'hb == _GEN_79 ? 1'h0 : registerTagMap_11_valid; // @[ReorderBuffer.scala 97:{13,13} 69:39]
  wire  _GEN_156 = 5'hc == _GEN_79 ? 1'h0 : registerTagMap_12_valid; // @[ReorderBuffer.scala 97:{13,13} 69:39]
  wire  _GEN_157 = 5'hd == _GEN_79 ? 1'h0 : registerTagMap_13_valid; // @[ReorderBuffer.scala 97:{13,13} 69:39]
  wire  _GEN_158 = 5'he == _GEN_79 ? 1'h0 : registerTagMap_14_valid; // @[ReorderBuffer.scala 97:{13,13} 69:39]
  wire  _GEN_159 = 5'hf == _GEN_79 ? 1'h0 : registerTagMap_15_valid; // @[ReorderBuffer.scala 97:{13,13} 69:39]
  wire  _GEN_160 = 5'h10 == _GEN_79 ? 1'h0 : registerTagMap_16_valid; // @[ReorderBuffer.scala 97:{13,13} 69:39]
  wire  _GEN_161 = 5'h11 == _GEN_79 ? 1'h0 : registerTagMap_17_valid; // @[ReorderBuffer.scala 97:{13,13} 69:39]
  wire  _GEN_162 = 5'h12 == _GEN_79 ? 1'h0 : registerTagMap_18_valid; // @[ReorderBuffer.scala 97:{13,13} 69:39]
  wire  _GEN_163 = 5'h13 == _GEN_79 ? 1'h0 : registerTagMap_19_valid; // @[ReorderBuffer.scala 97:{13,13} 69:39]
  wire  _GEN_164 = 5'h14 == _GEN_79 ? 1'h0 : registerTagMap_20_valid; // @[ReorderBuffer.scala 97:{13,13} 69:39]
  wire  _GEN_165 = 5'h15 == _GEN_79 ? 1'h0 : registerTagMap_21_valid; // @[ReorderBuffer.scala 97:{13,13} 69:39]
  wire  _GEN_166 = 5'h16 == _GEN_79 ? 1'h0 : registerTagMap_22_valid; // @[ReorderBuffer.scala 97:{13,13} 69:39]
  wire  _GEN_167 = 5'h17 == _GEN_79 ? 1'h0 : registerTagMap_23_valid; // @[ReorderBuffer.scala 97:{13,13} 69:39]
  wire  _GEN_168 = 5'h18 == _GEN_79 ? 1'h0 : registerTagMap_24_valid; // @[ReorderBuffer.scala 97:{13,13} 69:39]
  wire  _GEN_169 = 5'h19 == _GEN_79 ? 1'h0 : registerTagMap_25_valid; // @[ReorderBuffer.scala 97:{13,13} 69:39]
  wire  _GEN_170 = 5'h1a == _GEN_79 ? 1'h0 : registerTagMap_26_valid; // @[ReorderBuffer.scala 97:{13,13} 69:39]
  wire  _GEN_171 = 5'h1b == _GEN_79 ? 1'h0 : registerTagMap_27_valid; // @[ReorderBuffer.scala 97:{13,13} 69:39]
  wire  _GEN_172 = 5'h1c == _GEN_79 ? 1'h0 : registerTagMap_28_valid; // @[ReorderBuffer.scala 97:{13,13} 69:39]
  wire  _GEN_173 = 5'h1d == _GEN_79 ? 1'h0 : registerTagMap_29_valid; // @[ReorderBuffer.scala 97:{13,13} 69:39]
  wire  _GEN_174 = 5'h1e == _GEN_79 ? 1'h0 : registerTagMap_30_valid; // @[ReorderBuffer.scala 97:{13,13} 69:39]
  wire  _GEN_175 = 5'h1f == _GEN_79 ? 1'h0 : registerTagMap_31_valid; // @[ReorderBuffer.scala 97:{13,13} 69:39]
  wire  _GEN_177 = _T_1 ? _GEN_145 : registerTagMap_1_valid; // @[ReorderBuffer.scala 94:11 69:39]
  wire  _GEN_178 = _T_1 ? _GEN_146 : registerTagMap_2_valid; // @[ReorderBuffer.scala 94:11 69:39]
  wire  _GEN_179 = _T_1 ? _GEN_147 : registerTagMap_3_valid; // @[ReorderBuffer.scala 94:11 69:39]
  wire  _GEN_180 = _T_1 ? _GEN_148 : registerTagMap_4_valid; // @[ReorderBuffer.scala 94:11 69:39]
  wire  _GEN_181 = _T_1 ? _GEN_149 : registerTagMap_5_valid; // @[ReorderBuffer.scala 94:11 69:39]
  wire  _GEN_182 = _T_1 ? _GEN_150 : registerTagMap_6_valid; // @[ReorderBuffer.scala 94:11 69:39]
  wire  _GEN_183 = _T_1 ? _GEN_151 : registerTagMap_7_valid; // @[ReorderBuffer.scala 94:11 69:39]
  wire  _GEN_184 = _T_1 ? _GEN_152 : registerTagMap_8_valid; // @[ReorderBuffer.scala 94:11 69:39]
  wire  _GEN_185 = _T_1 ? _GEN_153 : registerTagMap_9_valid; // @[ReorderBuffer.scala 94:11 69:39]
  wire  _GEN_186 = _T_1 ? _GEN_154 : registerTagMap_10_valid; // @[ReorderBuffer.scala 94:11 69:39]
  wire  _GEN_187 = _T_1 ? _GEN_155 : registerTagMap_11_valid; // @[ReorderBuffer.scala 94:11 69:39]
  wire  _GEN_188 = _T_1 ? _GEN_156 : registerTagMap_12_valid; // @[ReorderBuffer.scala 94:11 69:39]
  wire  _GEN_189 = _T_1 ? _GEN_157 : registerTagMap_13_valid; // @[ReorderBuffer.scala 94:11 69:39]
  wire  _GEN_190 = _T_1 ? _GEN_158 : registerTagMap_14_valid; // @[ReorderBuffer.scala 94:11 69:39]
  wire  _GEN_191 = _T_1 ? _GEN_159 : registerTagMap_15_valid; // @[ReorderBuffer.scala 94:11 69:39]
  wire  _GEN_192 = _T_1 ? _GEN_160 : registerTagMap_16_valid; // @[ReorderBuffer.scala 94:11 69:39]
  wire  _GEN_193 = _T_1 ? _GEN_161 : registerTagMap_17_valid; // @[ReorderBuffer.scala 94:11 69:39]
  wire  _GEN_194 = _T_1 ? _GEN_162 : registerTagMap_18_valid; // @[ReorderBuffer.scala 94:11 69:39]
  wire  _GEN_195 = _T_1 ? _GEN_163 : registerTagMap_19_valid; // @[ReorderBuffer.scala 94:11 69:39]
  wire  _GEN_196 = _T_1 ? _GEN_164 : registerTagMap_20_valid; // @[ReorderBuffer.scala 94:11 69:39]
  wire  _GEN_197 = _T_1 ? _GEN_165 : registerTagMap_21_valid; // @[ReorderBuffer.scala 94:11 69:39]
  wire  _GEN_198 = _T_1 ? _GEN_166 : registerTagMap_22_valid; // @[ReorderBuffer.scala 94:11 69:39]
  wire  _GEN_199 = _T_1 ? _GEN_167 : registerTagMap_23_valid; // @[ReorderBuffer.scala 94:11 69:39]
  wire  _GEN_200 = _T_1 ? _GEN_168 : registerTagMap_24_valid; // @[ReorderBuffer.scala 94:11 69:39]
  wire  _GEN_201 = _T_1 ? _GEN_169 : registerTagMap_25_valid; // @[ReorderBuffer.scala 94:11 69:39]
  wire  _GEN_202 = _T_1 ? _GEN_170 : registerTagMap_26_valid; // @[ReorderBuffer.scala 94:11 69:39]
  wire  _GEN_203 = _T_1 ? _GEN_171 : registerTagMap_27_valid; // @[ReorderBuffer.scala 94:11 69:39]
  wire  _GEN_204 = _T_1 ? _GEN_172 : registerTagMap_28_valid; // @[ReorderBuffer.scala 94:11 69:39]
  wire  _GEN_205 = _T_1 ? _GEN_173 : registerTagMap_29_valid; // @[ReorderBuffer.scala 94:11 69:39]
  wire  _GEN_206 = _T_1 ? _GEN_174 : registerTagMap_30_valid; // @[ReorderBuffer.scala 94:11 69:39]
  wire  _GEN_207 = _T_1 ? _GEN_175 : registerTagMap_31_valid; // @[ReorderBuffer.scala 94:11 69:39]
  wire [63:0] _GEN_208 = _io_registerFile_0_valid_T ? _GEN_63 : 64'h0; // @[ReorderBuffer.scala 84:19 89:22 90:23]
  wire [4:0] _GEN_209 = _io_registerFile_0_valid_T ? _GEN_79 : 5'h0; // @[ReorderBuffer.scala 89:22 85:33 91:37]
  wire  _GEN_211 = _io_registerFile_0_valid_T ? _GEN_177 : registerTagMap_1_valid; // @[ReorderBuffer.scala 89:22 69:39]
  wire  _GEN_212 = _io_registerFile_0_valid_T ? _GEN_178 : registerTagMap_2_valid; // @[ReorderBuffer.scala 89:22 69:39]
  wire  _GEN_213 = _io_registerFile_0_valid_T ? _GEN_179 : registerTagMap_3_valid; // @[ReorderBuffer.scala 89:22 69:39]
  wire  _GEN_214 = _io_registerFile_0_valid_T ? _GEN_180 : registerTagMap_4_valid; // @[ReorderBuffer.scala 89:22 69:39]
  wire  _GEN_215 = _io_registerFile_0_valid_T ? _GEN_181 : registerTagMap_5_valid; // @[ReorderBuffer.scala 89:22 69:39]
  wire  _GEN_216 = _io_registerFile_0_valid_T ? _GEN_182 : registerTagMap_6_valid; // @[ReorderBuffer.scala 89:22 69:39]
  wire  _GEN_217 = _io_registerFile_0_valid_T ? _GEN_183 : registerTagMap_7_valid; // @[ReorderBuffer.scala 89:22 69:39]
  wire  _GEN_218 = _io_registerFile_0_valid_T ? _GEN_184 : registerTagMap_8_valid; // @[ReorderBuffer.scala 89:22 69:39]
  wire  _GEN_219 = _io_registerFile_0_valid_T ? _GEN_185 : registerTagMap_9_valid; // @[ReorderBuffer.scala 89:22 69:39]
  wire  _GEN_220 = _io_registerFile_0_valid_T ? _GEN_186 : registerTagMap_10_valid; // @[ReorderBuffer.scala 89:22 69:39]
  wire  _GEN_221 = _io_registerFile_0_valid_T ? _GEN_187 : registerTagMap_11_valid; // @[ReorderBuffer.scala 89:22 69:39]
  wire  _GEN_222 = _io_registerFile_0_valid_T ? _GEN_188 : registerTagMap_12_valid; // @[ReorderBuffer.scala 89:22 69:39]
  wire  _GEN_223 = _io_registerFile_0_valid_T ? _GEN_189 : registerTagMap_13_valid; // @[ReorderBuffer.scala 89:22 69:39]
  wire  _GEN_224 = _io_registerFile_0_valid_T ? _GEN_190 : registerTagMap_14_valid; // @[ReorderBuffer.scala 89:22 69:39]
  wire  _GEN_225 = _io_registerFile_0_valid_T ? _GEN_191 : registerTagMap_15_valid; // @[ReorderBuffer.scala 89:22 69:39]
  wire  _GEN_226 = _io_registerFile_0_valid_T ? _GEN_192 : registerTagMap_16_valid; // @[ReorderBuffer.scala 89:22 69:39]
  wire  _GEN_227 = _io_registerFile_0_valid_T ? _GEN_193 : registerTagMap_17_valid; // @[ReorderBuffer.scala 89:22 69:39]
  wire  _GEN_228 = _io_registerFile_0_valid_T ? _GEN_194 : registerTagMap_18_valid; // @[ReorderBuffer.scala 89:22 69:39]
  wire  _GEN_229 = _io_registerFile_0_valid_T ? _GEN_195 : registerTagMap_19_valid; // @[ReorderBuffer.scala 89:22 69:39]
  wire  _GEN_230 = _io_registerFile_0_valid_T ? _GEN_196 : registerTagMap_20_valid; // @[ReorderBuffer.scala 89:22 69:39]
  wire  _GEN_231 = _io_registerFile_0_valid_T ? _GEN_197 : registerTagMap_21_valid; // @[ReorderBuffer.scala 89:22 69:39]
  wire  _GEN_232 = _io_registerFile_0_valid_T ? _GEN_198 : registerTagMap_22_valid; // @[ReorderBuffer.scala 89:22 69:39]
  wire  _GEN_233 = _io_registerFile_0_valid_T ? _GEN_199 : registerTagMap_23_valid; // @[ReorderBuffer.scala 89:22 69:39]
  wire  _GEN_234 = _io_registerFile_0_valid_T ? _GEN_200 : registerTagMap_24_valid; // @[ReorderBuffer.scala 89:22 69:39]
  wire  _GEN_235 = _io_registerFile_0_valid_T ? _GEN_201 : registerTagMap_25_valid; // @[ReorderBuffer.scala 89:22 69:39]
  wire  _GEN_236 = _io_registerFile_0_valid_T ? _GEN_202 : registerTagMap_26_valid; // @[ReorderBuffer.scala 89:22 69:39]
  wire  _GEN_237 = _io_registerFile_0_valid_T ? _GEN_203 : registerTagMap_27_valid; // @[ReorderBuffer.scala 89:22 69:39]
  wire  _GEN_238 = _io_registerFile_0_valid_T ? _GEN_204 : registerTagMap_28_valid; // @[ReorderBuffer.scala 89:22 69:39]
  wire  _GEN_239 = _io_registerFile_0_valid_T ? _GEN_205 : registerTagMap_29_valid; // @[ReorderBuffer.scala 89:22 69:39]
  wire  _GEN_240 = _io_registerFile_0_valid_T ? _GEN_206 : registerTagMap_30_valid; // @[ReorderBuffer.scala 89:22 69:39]
  wire  _GEN_241 = _io_registerFile_0_valid_T ? _GEN_207 : registerTagMap_31_valid; // @[ReorderBuffer.scala 89:22 69:39]
  wire  _GEN_242 = _io_registerFile_0_valid_T ? 1'h0 : 1'h1; // @[ReorderBuffer.scala 89:22 86:25 100:29]
  wire  _GEN_247 = canCommit ? _GEN_211 : registerTagMap_1_valid; // @[ReorderBuffer.scala 88:21 69:39]
  wire  _GEN_248 = canCommit ? _GEN_212 : registerTagMap_2_valid; // @[ReorderBuffer.scala 88:21 69:39]
  wire  _GEN_249 = canCommit ? _GEN_213 : registerTagMap_3_valid; // @[ReorderBuffer.scala 88:21 69:39]
  wire  _GEN_250 = canCommit ? _GEN_214 : registerTagMap_4_valid; // @[ReorderBuffer.scala 88:21 69:39]
  wire  _GEN_251 = canCommit ? _GEN_215 : registerTagMap_5_valid; // @[ReorderBuffer.scala 88:21 69:39]
  wire  _GEN_252 = canCommit ? _GEN_216 : registerTagMap_6_valid; // @[ReorderBuffer.scala 88:21 69:39]
  wire  _GEN_253 = canCommit ? _GEN_217 : registerTagMap_7_valid; // @[ReorderBuffer.scala 88:21 69:39]
  wire  _GEN_254 = canCommit ? _GEN_218 : registerTagMap_8_valid; // @[ReorderBuffer.scala 88:21 69:39]
  wire  _GEN_255 = canCommit ? _GEN_219 : registerTagMap_9_valid; // @[ReorderBuffer.scala 88:21 69:39]
  wire  _GEN_256 = canCommit ? _GEN_220 : registerTagMap_10_valid; // @[ReorderBuffer.scala 88:21 69:39]
  wire  _GEN_257 = canCommit ? _GEN_221 : registerTagMap_11_valid; // @[ReorderBuffer.scala 88:21 69:39]
  wire  _GEN_258 = canCommit ? _GEN_222 : registerTagMap_12_valid; // @[ReorderBuffer.scala 88:21 69:39]
  wire  _GEN_259 = canCommit ? _GEN_223 : registerTagMap_13_valid; // @[ReorderBuffer.scala 88:21 69:39]
  wire  _GEN_260 = canCommit ? _GEN_224 : registerTagMap_14_valid; // @[ReorderBuffer.scala 88:21 69:39]
  wire  _GEN_261 = canCommit ? _GEN_225 : registerTagMap_15_valid; // @[ReorderBuffer.scala 88:21 69:39]
  wire  _GEN_262 = canCommit ? _GEN_226 : registerTagMap_16_valid; // @[ReorderBuffer.scala 88:21 69:39]
  wire  _GEN_263 = canCommit ? _GEN_227 : registerTagMap_17_valid; // @[ReorderBuffer.scala 88:21 69:39]
  wire  _GEN_264 = canCommit ? _GEN_228 : registerTagMap_18_valid; // @[ReorderBuffer.scala 88:21 69:39]
  wire  _GEN_265 = canCommit ? _GEN_229 : registerTagMap_19_valid; // @[ReorderBuffer.scala 88:21 69:39]
  wire  _GEN_266 = canCommit ? _GEN_230 : registerTagMap_20_valid; // @[ReorderBuffer.scala 88:21 69:39]
  wire  _GEN_267 = canCommit ? _GEN_231 : registerTagMap_21_valid; // @[ReorderBuffer.scala 88:21 69:39]
  wire  _GEN_268 = canCommit ? _GEN_232 : registerTagMap_22_valid; // @[ReorderBuffer.scala 88:21 69:39]
  wire  _GEN_269 = canCommit ? _GEN_233 : registerTagMap_23_valid; // @[ReorderBuffer.scala 88:21 69:39]
  wire  _GEN_270 = canCommit ? _GEN_234 : registerTagMap_24_valid; // @[ReorderBuffer.scala 88:21 69:39]
  wire  _GEN_271 = canCommit ? _GEN_235 : registerTagMap_25_valid; // @[ReorderBuffer.scala 88:21 69:39]
  wire  _GEN_272 = canCommit ? _GEN_236 : registerTagMap_26_valid; // @[ReorderBuffer.scala 88:21 69:39]
  wire  _GEN_273 = canCommit ? _GEN_237 : registerTagMap_27_valid; // @[ReorderBuffer.scala 88:21 69:39]
  wire  _GEN_274 = canCommit ? _GEN_238 : registerTagMap_28_valid; // @[ReorderBuffer.scala 88:21 69:39]
  wire  _GEN_275 = canCommit ? _GEN_239 : registerTagMap_29_valid; // @[ReorderBuffer.scala 88:21 69:39]
  wire  _GEN_276 = canCommit ? _GEN_240 : registerTagMap_30_valid; // @[ReorderBuffer.scala 88:21 69:39]
  wire  _GEN_277 = canCommit ? _GEN_241 : registerTagMap_31_valid; // @[ReorderBuffer.scala 88:21 69:39]
  wire  _GEN_278 = canCommit & _GEN_242; // @[ReorderBuffer.scala 88:21 86:25]
  wire [3:0] index_1 = tail + 4'h1; // @[ReorderBuffer.scala 77:22]
  wire  _GEN_300 = 4'h1 == index_1 ? buffer_1_valueReady : buffer_0_valueReady; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_301 = 4'h2 == index_1 ? buffer_2_valueReady : _GEN_300; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_302 = 4'h3 == index_1 ? buffer_3_valueReady : _GEN_301; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_303 = 4'h4 == index_1 ? buffer_4_valueReady : _GEN_302; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_304 = 4'h5 == index_1 ? buffer_5_valueReady : _GEN_303; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_305 = 4'h6 == index_1 ? buffer_6_valueReady : _GEN_304; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_306 = 4'h7 == index_1 ? buffer_7_valueReady : _GEN_305; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_307 = 4'h8 == index_1 ? buffer_8_valueReady : _GEN_306; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_308 = 4'h9 == index_1 ? buffer_9_valueReady : _GEN_307; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_309 = 4'ha == index_1 ? buffer_10_valueReady : _GEN_308; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_310 = 4'hb == index_1 ? buffer_11_valueReady : _GEN_309; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_311 = 4'hc == index_1 ? buffer_12_valueReady : _GEN_310; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_312 = 4'hd == index_1 ? buffer_13_valueReady : _GEN_311; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_313 = 4'he == index_1 ? buffer_14_valueReady : _GEN_312; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_314 = 4'hf == index_1 ? buffer_15_valueReady : _GEN_313; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_316 = 4'h1 == index_1 ? buffer_1_storeSign : buffer_0_storeSign; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_317 = 4'h2 == index_1 ? buffer_2_storeSign : _GEN_316; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_318 = 4'h3 == index_1 ? buffer_3_storeSign : _GEN_317; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_319 = 4'h4 == index_1 ? buffer_4_storeSign : _GEN_318; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_320 = 4'h5 == index_1 ? buffer_5_storeSign : _GEN_319; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_321 = 4'h6 == index_1 ? buffer_6_storeSign : _GEN_320; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_322 = 4'h7 == index_1 ? buffer_7_storeSign : _GEN_321; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_323 = 4'h8 == index_1 ? buffer_8_storeSign : _GEN_322; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_324 = 4'h9 == index_1 ? buffer_9_storeSign : _GEN_323; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_325 = 4'ha == index_1 ? buffer_10_storeSign : _GEN_324; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_326 = 4'hb == index_1 ? buffer_11_storeSign : _GEN_325; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_327 = 4'hc == index_1 ? buffer_12_storeSign : _GEN_326; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_328 = 4'hd == index_1 ? buffer_13_storeSign : _GEN_327; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_329 = 4'he == index_1 ? buffer_14_storeSign : _GEN_328; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_330 = 4'hf == index_1 ? buffer_15_storeSign : _GEN_329; // @[ReorderBuffer.scala 79:{50,50}]
  wire  instructionOk_1 = _GEN_314 | _GEN_330; // @[ReorderBuffer.scala 79:50]
  wire  canCommit_1 = canCommit & index_1 != head & instructionOk_1; // @[ReorderBuffer.scala 80:49]
  wire  _GEN_332 = 4'h1 == index_1 ? buffer_1_isError : buffer_0_isError; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_333 = 4'h2 == index_1 ? buffer_2_isError : _GEN_332; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_334 = 4'h3 == index_1 ? buffer_3_isError : _GEN_333; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_335 = 4'h4 == index_1 ? buffer_4_isError : _GEN_334; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_336 = 4'h5 == index_1 ? buffer_5_isError : _GEN_335; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_337 = 4'h6 == index_1 ? buffer_6_isError : _GEN_336; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_338 = 4'h7 == index_1 ? buffer_7_isError : _GEN_337; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_339 = 4'h8 == index_1 ? buffer_8_isError : _GEN_338; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_340 = 4'h9 == index_1 ? buffer_9_isError : _GEN_339; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_341 = 4'ha == index_1 ? buffer_10_isError : _GEN_340; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_342 = 4'hb == index_1 ? buffer_11_isError : _GEN_341; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_343 = 4'hc == index_1 ? buffer_12_isError : _GEN_342; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_344 = 4'hd == index_1 ? buffer_13_isError : _GEN_343; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_345 = 4'he == index_1 ? buffer_14_isError : _GEN_344; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_346 = 4'hf == index_1 ? buffer_15_isError : _GEN_345; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _io_registerFile_1_valid_T = ~_GEN_346; // @[ReorderBuffer.scala 83:30]
  wire [63:0] _GEN_348 = 4'h1 == index_1 ? buffer_1_value : buffer_0_value; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_349 = 4'h2 == index_1 ? buffer_2_value : _GEN_348; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_350 = 4'h3 == index_1 ? buffer_3_value : _GEN_349; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_351 = 4'h4 == index_1 ? buffer_4_value : _GEN_350; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_352 = 4'h5 == index_1 ? buffer_5_value : _GEN_351; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_353 = 4'h6 == index_1 ? buffer_6_value : _GEN_352; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_354 = 4'h7 == index_1 ? buffer_7_value : _GEN_353; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_355 = 4'h8 == index_1 ? buffer_8_value : _GEN_354; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_356 = 4'h9 == index_1 ? buffer_9_value : _GEN_355; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_357 = 4'ha == index_1 ? buffer_10_value : _GEN_356; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_358 = 4'hb == index_1 ? buffer_11_value : _GEN_357; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_359 = 4'hc == index_1 ? buffer_12_value : _GEN_358; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_360 = 4'hd == index_1 ? buffer_13_value : _GEN_359; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_361 = 4'he == index_1 ? buffer_14_value : _GEN_360; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_362 = 4'hf == index_1 ? buffer_15_value : _GEN_361; // @[ReorderBuffer.scala 90:{23,23}]
  wire [4:0] _GEN_364 = 4'h1 == index_1 ? buffer_1_destinationRegister : buffer_0_destinationRegister; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_365 = 4'h2 == index_1 ? buffer_2_destinationRegister : _GEN_364; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_366 = 4'h3 == index_1 ? buffer_3_destinationRegister : _GEN_365; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_367 = 4'h4 == index_1 ? buffer_4_destinationRegister : _GEN_366; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_368 = 4'h5 == index_1 ? buffer_5_destinationRegister : _GEN_367; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_369 = 4'h6 == index_1 ? buffer_6_destinationRegister : _GEN_368; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_370 = 4'h7 == index_1 ? buffer_7_destinationRegister : _GEN_369; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_371 = 4'h8 == index_1 ? buffer_8_destinationRegister : _GEN_370; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_372 = 4'h9 == index_1 ? buffer_9_destinationRegister : _GEN_371; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_373 = 4'ha == index_1 ? buffer_10_destinationRegister : _GEN_372; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_374 = 4'hb == index_1 ? buffer_11_destinationRegister : _GEN_373; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_375 = 4'hc == index_1 ? buffer_12_destinationRegister : _GEN_374; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_376 = 4'hd == index_1 ? buffer_13_destinationRegister : _GEN_375; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_377 = 4'he == index_1 ? buffer_14_destinationRegister : _GEN_376; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_378 = 4'hf == index_1 ? buffer_15_destinationRegister : _GEN_377; // @[ReorderBuffer.scala 91:{37,37}]
  wire [3:0] _GEN_380 = 5'h1 == _GEN_378 ? registerTagMap_1_tagId : 4'h0; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_381 = 5'h2 == _GEN_378 ? registerTagMap_2_tagId : _GEN_380; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_382 = 5'h3 == _GEN_378 ? registerTagMap_3_tagId : _GEN_381; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_383 = 5'h4 == _GEN_378 ? registerTagMap_4_tagId : _GEN_382; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_384 = 5'h5 == _GEN_378 ? registerTagMap_5_tagId : _GEN_383; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_385 = 5'h6 == _GEN_378 ? registerTagMap_6_tagId : _GEN_384; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_386 = 5'h7 == _GEN_378 ? registerTagMap_7_tagId : _GEN_385; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_387 = 5'h8 == _GEN_378 ? registerTagMap_8_tagId : _GEN_386; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_388 = 5'h9 == _GEN_378 ? registerTagMap_9_tagId : _GEN_387; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_389 = 5'ha == _GEN_378 ? registerTagMap_10_tagId : _GEN_388; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_390 = 5'hb == _GEN_378 ? registerTagMap_11_tagId : _GEN_389; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_391 = 5'hc == _GEN_378 ? registerTagMap_12_tagId : _GEN_390; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_392 = 5'hd == _GEN_378 ? registerTagMap_13_tagId : _GEN_391; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_393 = 5'he == _GEN_378 ? registerTagMap_14_tagId : _GEN_392; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_394 = 5'hf == _GEN_378 ? registerTagMap_15_tagId : _GEN_393; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_395 = 5'h10 == _GEN_378 ? registerTagMap_16_tagId : _GEN_394; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_396 = 5'h11 == _GEN_378 ? registerTagMap_17_tagId : _GEN_395; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_397 = 5'h12 == _GEN_378 ? registerTagMap_18_tagId : _GEN_396; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_398 = 5'h13 == _GEN_378 ? registerTagMap_19_tagId : _GEN_397; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_399 = 5'h14 == _GEN_378 ? registerTagMap_20_tagId : _GEN_398; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_400 = 5'h15 == _GEN_378 ? registerTagMap_21_tagId : _GEN_399; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_401 = 5'h16 == _GEN_378 ? registerTagMap_22_tagId : _GEN_400; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_402 = 5'h17 == _GEN_378 ? registerTagMap_23_tagId : _GEN_401; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_403 = 5'h18 == _GEN_378 ? registerTagMap_24_tagId : _GEN_402; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_404 = 5'h19 == _GEN_378 ? registerTagMap_25_tagId : _GEN_403; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_405 = 5'h1a == _GEN_378 ? registerTagMap_26_tagId : _GEN_404; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_406 = 5'h1b == _GEN_378 ? registerTagMap_27_tagId : _GEN_405; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_407 = 5'h1c == _GEN_378 ? registerTagMap_28_tagId : _GEN_406; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_408 = 5'h1d == _GEN_378 ? registerTagMap_29_tagId : _GEN_407; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_409 = 5'h1e == _GEN_378 ? registerTagMap_30_tagId : _GEN_408; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_410 = 5'h1f == _GEN_378 ? registerTagMap_31_tagId : _GEN_409; // @[ReorderBuffer.scala 93:{17,17}]
  wire  _T_3 = index_1 == _GEN_410; // @[ReorderBuffer.scala 93:17]
  wire  _GEN_444 = 5'h1 == _GEN_378 ? 1'h0 : _GEN_247; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_445 = 5'h2 == _GEN_378 ? 1'h0 : _GEN_248; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_446 = 5'h3 == _GEN_378 ? 1'h0 : _GEN_249; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_447 = 5'h4 == _GEN_378 ? 1'h0 : _GEN_250; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_448 = 5'h5 == _GEN_378 ? 1'h0 : _GEN_251; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_449 = 5'h6 == _GEN_378 ? 1'h0 : _GEN_252; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_450 = 5'h7 == _GEN_378 ? 1'h0 : _GEN_253; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_451 = 5'h8 == _GEN_378 ? 1'h0 : _GEN_254; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_452 = 5'h9 == _GEN_378 ? 1'h0 : _GEN_255; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_453 = 5'ha == _GEN_378 ? 1'h0 : _GEN_256; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_454 = 5'hb == _GEN_378 ? 1'h0 : _GEN_257; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_455 = 5'hc == _GEN_378 ? 1'h0 : _GEN_258; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_456 = 5'hd == _GEN_378 ? 1'h0 : _GEN_259; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_457 = 5'he == _GEN_378 ? 1'h0 : _GEN_260; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_458 = 5'hf == _GEN_378 ? 1'h0 : _GEN_261; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_459 = 5'h10 == _GEN_378 ? 1'h0 : _GEN_262; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_460 = 5'h11 == _GEN_378 ? 1'h0 : _GEN_263; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_461 = 5'h12 == _GEN_378 ? 1'h0 : _GEN_264; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_462 = 5'h13 == _GEN_378 ? 1'h0 : _GEN_265; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_463 = 5'h14 == _GEN_378 ? 1'h0 : _GEN_266; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_464 = 5'h15 == _GEN_378 ? 1'h0 : _GEN_267; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_465 = 5'h16 == _GEN_378 ? 1'h0 : _GEN_268; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_466 = 5'h17 == _GEN_378 ? 1'h0 : _GEN_269; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_467 = 5'h18 == _GEN_378 ? 1'h0 : _GEN_270; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_468 = 5'h19 == _GEN_378 ? 1'h0 : _GEN_271; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_469 = 5'h1a == _GEN_378 ? 1'h0 : _GEN_272; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_470 = 5'h1b == _GEN_378 ? 1'h0 : _GEN_273; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_471 = 5'h1c == _GEN_378 ? 1'h0 : _GEN_274; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_472 = 5'h1d == _GEN_378 ? 1'h0 : _GEN_275; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_473 = 5'h1e == _GEN_378 ? 1'h0 : _GEN_276; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_474 = 5'h1f == _GEN_378 ? 1'h0 : _GEN_277; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_476 = _T_3 ? _GEN_444 : _GEN_247; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_477 = _T_3 ? _GEN_445 : _GEN_248; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_478 = _T_3 ? _GEN_446 : _GEN_249; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_479 = _T_3 ? _GEN_447 : _GEN_250; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_480 = _T_3 ? _GEN_448 : _GEN_251; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_481 = _T_3 ? _GEN_449 : _GEN_252; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_482 = _T_3 ? _GEN_450 : _GEN_253; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_483 = _T_3 ? _GEN_451 : _GEN_254; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_484 = _T_3 ? _GEN_452 : _GEN_255; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_485 = _T_3 ? _GEN_453 : _GEN_256; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_486 = _T_3 ? _GEN_454 : _GEN_257; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_487 = _T_3 ? _GEN_455 : _GEN_258; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_488 = _T_3 ? _GEN_456 : _GEN_259; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_489 = _T_3 ? _GEN_457 : _GEN_260; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_490 = _T_3 ? _GEN_458 : _GEN_261; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_491 = _T_3 ? _GEN_459 : _GEN_262; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_492 = _T_3 ? _GEN_460 : _GEN_263; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_493 = _T_3 ? _GEN_461 : _GEN_264; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_494 = _T_3 ? _GEN_462 : _GEN_265; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_495 = _T_3 ? _GEN_463 : _GEN_266; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_496 = _T_3 ? _GEN_464 : _GEN_267; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_497 = _T_3 ? _GEN_465 : _GEN_268; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_498 = _T_3 ? _GEN_466 : _GEN_269; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_499 = _T_3 ? _GEN_467 : _GEN_270; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_500 = _T_3 ? _GEN_468 : _GEN_271; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_501 = _T_3 ? _GEN_469 : _GEN_272; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_502 = _T_3 ? _GEN_470 : _GEN_273; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_503 = _T_3 ? _GEN_471 : _GEN_274; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_504 = _T_3 ? _GEN_472 : _GEN_275; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_505 = _T_3 ? _GEN_473 : _GEN_276; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_506 = _T_3 ? _GEN_474 : _GEN_277; // @[ReorderBuffer.scala 94:11]
  wire [63:0] _GEN_507 = _io_registerFile_1_valid_T ? _GEN_362 : 64'h0; // @[ReorderBuffer.scala 84:19 89:22 90:23]
  wire [4:0] _GEN_508 = _io_registerFile_1_valid_T ? _GEN_378 : 5'h0; // @[ReorderBuffer.scala 89:22 85:33 91:37]
  wire  _GEN_510 = _io_registerFile_1_valid_T ? _GEN_476 : _GEN_247; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_511 = _io_registerFile_1_valid_T ? _GEN_477 : _GEN_248; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_512 = _io_registerFile_1_valid_T ? _GEN_478 : _GEN_249; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_513 = _io_registerFile_1_valid_T ? _GEN_479 : _GEN_250; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_514 = _io_registerFile_1_valid_T ? _GEN_480 : _GEN_251; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_515 = _io_registerFile_1_valid_T ? _GEN_481 : _GEN_252; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_516 = _io_registerFile_1_valid_T ? _GEN_482 : _GEN_253; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_517 = _io_registerFile_1_valid_T ? _GEN_483 : _GEN_254; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_518 = _io_registerFile_1_valid_T ? _GEN_484 : _GEN_255; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_519 = _io_registerFile_1_valid_T ? _GEN_485 : _GEN_256; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_520 = _io_registerFile_1_valid_T ? _GEN_486 : _GEN_257; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_521 = _io_registerFile_1_valid_T ? _GEN_487 : _GEN_258; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_522 = _io_registerFile_1_valid_T ? _GEN_488 : _GEN_259; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_523 = _io_registerFile_1_valid_T ? _GEN_489 : _GEN_260; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_524 = _io_registerFile_1_valid_T ? _GEN_490 : _GEN_261; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_525 = _io_registerFile_1_valid_T ? _GEN_491 : _GEN_262; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_526 = _io_registerFile_1_valid_T ? _GEN_492 : _GEN_263; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_527 = _io_registerFile_1_valid_T ? _GEN_493 : _GEN_264; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_528 = _io_registerFile_1_valid_T ? _GEN_494 : _GEN_265; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_529 = _io_registerFile_1_valid_T ? _GEN_495 : _GEN_266; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_530 = _io_registerFile_1_valid_T ? _GEN_496 : _GEN_267; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_531 = _io_registerFile_1_valid_T ? _GEN_497 : _GEN_268; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_532 = _io_registerFile_1_valid_T ? _GEN_498 : _GEN_269; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_533 = _io_registerFile_1_valid_T ? _GEN_499 : _GEN_270; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_534 = _io_registerFile_1_valid_T ? _GEN_500 : _GEN_271; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_535 = _io_registerFile_1_valid_T ? _GEN_501 : _GEN_272; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_536 = _io_registerFile_1_valid_T ? _GEN_502 : _GEN_273; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_537 = _io_registerFile_1_valid_T ? _GEN_503 : _GEN_274; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_538 = _io_registerFile_1_valid_T ? _GEN_504 : _GEN_275; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_539 = _io_registerFile_1_valid_T ? _GEN_505 : _GEN_276; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_540 = _io_registerFile_1_valid_T ? _GEN_506 : _GEN_277; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_543 = _io_registerFile_1_valid_T ? _GEN_278 : 1'h1; // @[ReorderBuffer.scala 102:20 89:22]
  wire  _GEN_547 = canCommit_1 ? _GEN_510 : _GEN_247; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_548 = canCommit_1 ? _GEN_511 : _GEN_248; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_549 = canCommit_1 ? _GEN_512 : _GEN_249; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_550 = canCommit_1 ? _GEN_513 : _GEN_250; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_551 = canCommit_1 ? _GEN_514 : _GEN_251; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_552 = canCommit_1 ? _GEN_515 : _GEN_252; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_553 = canCommit_1 ? _GEN_516 : _GEN_253; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_554 = canCommit_1 ? _GEN_517 : _GEN_254; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_555 = canCommit_1 ? _GEN_518 : _GEN_255; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_556 = canCommit_1 ? _GEN_519 : _GEN_256; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_557 = canCommit_1 ? _GEN_520 : _GEN_257; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_558 = canCommit_1 ? _GEN_521 : _GEN_258; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_559 = canCommit_1 ? _GEN_522 : _GEN_259; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_560 = canCommit_1 ? _GEN_523 : _GEN_260; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_561 = canCommit_1 ? _GEN_524 : _GEN_261; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_562 = canCommit_1 ? _GEN_525 : _GEN_262; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_563 = canCommit_1 ? _GEN_526 : _GEN_263; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_564 = canCommit_1 ? _GEN_527 : _GEN_264; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_565 = canCommit_1 ? _GEN_528 : _GEN_265; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_566 = canCommit_1 ? _GEN_529 : _GEN_266; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_567 = canCommit_1 ? _GEN_530 : _GEN_267; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_568 = canCommit_1 ? _GEN_531 : _GEN_268; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_569 = canCommit_1 ? _GEN_532 : _GEN_269; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_570 = canCommit_1 ? _GEN_533 : _GEN_270; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_571 = canCommit_1 ? _GEN_534 : _GEN_271; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_572 = canCommit_1 ? _GEN_535 : _GEN_272; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_573 = canCommit_1 ? _GEN_536 : _GEN_273; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_574 = canCommit_1 ? _GEN_537 : _GEN_274; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_575 = canCommit_1 ? _GEN_538 : _GEN_275; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_576 = canCommit_1 ? _GEN_539 : _GEN_276; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_577 = canCommit_1 ? _GEN_540 : _GEN_277; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_580 = canCommit_1 ? _GEN_543 : _GEN_278; // @[ReorderBuffer.scala 88:21]
  wire [3:0] index_2 = tail + 4'h2; // @[ReorderBuffer.scala 77:22]
  wire  _GEN_601 = 4'h1 == index_2 ? buffer_1_valueReady : buffer_0_valueReady; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_602 = 4'h2 == index_2 ? buffer_2_valueReady : _GEN_601; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_603 = 4'h3 == index_2 ? buffer_3_valueReady : _GEN_602; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_604 = 4'h4 == index_2 ? buffer_4_valueReady : _GEN_603; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_605 = 4'h5 == index_2 ? buffer_5_valueReady : _GEN_604; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_606 = 4'h6 == index_2 ? buffer_6_valueReady : _GEN_605; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_607 = 4'h7 == index_2 ? buffer_7_valueReady : _GEN_606; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_608 = 4'h8 == index_2 ? buffer_8_valueReady : _GEN_607; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_609 = 4'h9 == index_2 ? buffer_9_valueReady : _GEN_608; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_610 = 4'ha == index_2 ? buffer_10_valueReady : _GEN_609; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_611 = 4'hb == index_2 ? buffer_11_valueReady : _GEN_610; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_612 = 4'hc == index_2 ? buffer_12_valueReady : _GEN_611; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_613 = 4'hd == index_2 ? buffer_13_valueReady : _GEN_612; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_614 = 4'he == index_2 ? buffer_14_valueReady : _GEN_613; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_615 = 4'hf == index_2 ? buffer_15_valueReady : _GEN_614; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_617 = 4'h1 == index_2 ? buffer_1_storeSign : buffer_0_storeSign; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_618 = 4'h2 == index_2 ? buffer_2_storeSign : _GEN_617; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_619 = 4'h3 == index_2 ? buffer_3_storeSign : _GEN_618; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_620 = 4'h4 == index_2 ? buffer_4_storeSign : _GEN_619; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_621 = 4'h5 == index_2 ? buffer_5_storeSign : _GEN_620; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_622 = 4'h6 == index_2 ? buffer_6_storeSign : _GEN_621; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_623 = 4'h7 == index_2 ? buffer_7_storeSign : _GEN_622; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_624 = 4'h8 == index_2 ? buffer_8_storeSign : _GEN_623; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_625 = 4'h9 == index_2 ? buffer_9_storeSign : _GEN_624; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_626 = 4'ha == index_2 ? buffer_10_storeSign : _GEN_625; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_627 = 4'hb == index_2 ? buffer_11_storeSign : _GEN_626; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_628 = 4'hc == index_2 ? buffer_12_storeSign : _GEN_627; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_629 = 4'hd == index_2 ? buffer_13_storeSign : _GEN_628; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_630 = 4'he == index_2 ? buffer_14_storeSign : _GEN_629; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_631 = 4'hf == index_2 ? buffer_15_storeSign : _GEN_630; // @[ReorderBuffer.scala 79:{50,50}]
  wire  instructionOk_2 = _GEN_615 | _GEN_631; // @[ReorderBuffer.scala 79:50]
  wire  canCommit_2 = canCommit_1 & index_2 != head & instructionOk_2; // @[ReorderBuffer.scala 80:49]
  wire  _GEN_633 = 4'h1 == index_2 ? buffer_1_isError : buffer_0_isError; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_634 = 4'h2 == index_2 ? buffer_2_isError : _GEN_633; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_635 = 4'h3 == index_2 ? buffer_3_isError : _GEN_634; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_636 = 4'h4 == index_2 ? buffer_4_isError : _GEN_635; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_637 = 4'h5 == index_2 ? buffer_5_isError : _GEN_636; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_638 = 4'h6 == index_2 ? buffer_6_isError : _GEN_637; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_639 = 4'h7 == index_2 ? buffer_7_isError : _GEN_638; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_640 = 4'h8 == index_2 ? buffer_8_isError : _GEN_639; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_641 = 4'h9 == index_2 ? buffer_9_isError : _GEN_640; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_642 = 4'ha == index_2 ? buffer_10_isError : _GEN_641; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_643 = 4'hb == index_2 ? buffer_11_isError : _GEN_642; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_644 = 4'hc == index_2 ? buffer_12_isError : _GEN_643; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_645 = 4'hd == index_2 ? buffer_13_isError : _GEN_644; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_646 = 4'he == index_2 ? buffer_14_isError : _GEN_645; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_647 = 4'hf == index_2 ? buffer_15_isError : _GEN_646; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _io_registerFile_2_valid_T = ~_GEN_647; // @[ReorderBuffer.scala 83:30]
  wire [63:0] _GEN_649 = 4'h1 == index_2 ? buffer_1_value : buffer_0_value; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_650 = 4'h2 == index_2 ? buffer_2_value : _GEN_649; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_651 = 4'h3 == index_2 ? buffer_3_value : _GEN_650; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_652 = 4'h4 == index_2 ? buffer_4_value : _GEN_651; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_653 = 4'h5 == index_2 ? buffer_5_value : _GEN_652; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_654 = 4'h6 == index_2 ? buffer_6_value : _GEN_653; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_655 = 4'h7 == index_2 ? buffer_7_value : _GEN_654; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_656 = 4'h8 == index_2 ? buffer_8_value : _GEN_655; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_657 = 4'h9 == index_2 ? buffer_9_value : _GEN_656; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_658 = 4'ha == index_2 ? buffer_10_value : _GEN_657; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_659 = 4'hb == index_2 ? buffer_11_value : _GEN_658; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_660 = 4'hc == index_2 ? buffer_12_value : _GEN_659; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_661 = 4'hd == index_2 ? buffer_13_value : _GEN_660; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_662 = 4'he == index_2 ? buffer_14_value : _GEN_661; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_663 = 4'hf == index_2 ? buffer_15_value : _GEN_662; // @[ReorderBuffer.scala 90:{23,23}]
  wire [4:0] _GEN_665 = 4'h1 == index_2 ? buffer_1_destinationRegister : buffer_0_destinationRegister; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_666 = 4'h2 == index_2 ? buffer_2_destinationRegister : _GEN_665; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_667 = 4'h3 == index_2 ? buffer_3_destinationRegister : _GEN_666; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_668 = 4'h4 == index_2 ? buffer_4_destinationRegister : _GEN_667; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_669 = 4'h5 == index_2 ? buffer_5_destinationRegister : _GEN_668; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_670 = 4'h6 == index_2 ? buffer_6_destinationRegister : _GEN_669; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_671 = 4'h7 == index_2 ? buffer_7_destinationRegister : _GEN_670; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_672 = 4'h8 == index_2 ? buffer_8_destinationRegister : _GEN_671; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_673 = 4'h9 == index_2 ? buffer_9_destinationRegister : _GEN_672; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_674 = 4'ha == index_2 ? buffer_10_destinationRegister : _GEN_673; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_675 = 4'hb == index_2 ? buffer_11_destinationRegister : _GEN_674; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_676 = 4'hc == index_2 ? buffer_12_destinationRegister : _GEN_675; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_677 = 4'hd == index_2 ? buffer_13_destinationRegister : _GEN_676; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_678 = 4'he == index_2 ? buffer_14_destinationRegister : _GEN_677; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_679 = 4'hf == index_2 ? buffer_15_destinationRegister : _GEN_678; // @[ReorderBuffer.scala 91:{37,37}]
  wire [3:0] _GEN_681 = 5'h1 == _GEN_679 ? registerTagMap_1_tagId : 4'h0; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_682 = 5'h2 == _GEN_679 ? registerTagMap_2_tagId : _GEN_681; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_683 = 5'h3 == _GEN_679 ? registerTagMap_3_tagId : _GEN_682; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_684 = 5'h4 == _GEN_679 ? registerTagMap_4_tagId : _GEN_683; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_685 = 5'h5 == _GEN_679 ? registerTagMap_5_tagId : _GEN_684; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_686 = 5'h6 == _GEN_679 ? registerTagMap_6_tagId : _GEN_685; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_687 = 5'h7 == _GEN_679 ? registerTagMap_7_tagId : _GEN_686; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_688 = 5'h8 == _GEN_679 ? registerTagMap_8_tagId : _GEN_687; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_689 = 5'h9 == _GEN_679 ? registerTagMap_9_tagId : _GEN_688; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_690 = 5'ha == _GEN_679 ? registerTagMap_10_tagId : _GEN_689; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_691 = 5'hb == _GEN_679 ? registerTagMap_11_tagId : _GEN_690; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_692 = 5'hc == _GEN_679 ? registerTagMap_12_tagId : _GEN_691; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_693 = 5'hd == _GEN_679 ? registerTagMap_13_tagId : _GEN_692; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_694 = 5'he == _GEN_679 ? registerTagMap_14_tagId : _GEN_693; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_695 = 5'hf == _GEN_679 ? registerTagMap_15_tagId : _GEN_694; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_696 = 5'h10 == _GEN_679 ? registerTagMap_16_tagId : _GEN_695; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_697 = 5'h11 == _GEN_679 ? registerTagMap_17_tagId : _GEN_696; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_698 = 5'h12 == _GEN_679 ? registerTagMap_18_tagId : _GEN_697; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_699 = 5'h13 == _GEN_679 ? registerTagMap_19_tagId : _GEN_698; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_700 = 5'h14 == _GEN_679 ? registerTagMap_20_tagId : _GEN_699; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_701 = 5'h15 == _GEN_679 ? registerTagMap_21_tagId : _GEN_700; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_702 = 5'h16 == _GEN_679 ? registerTagMap_22_tagId : _GEN_701; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_703 = 5'h17 == _GEN_679 ? registerTagMap_23_tagId : _GEN_702; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_704 = 5'h18 == _GEN_679 ? registerTagMap_24_tagId : _GEN_703; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_705 = 5'h19 == _GEN_679 ? registerTagMap_25_tagId : _GEN_704; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_706 = 5'h1a == _GEN_679 ? registerTagMap_26_tagId : _GEN_705; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_707 = 5'h1b == _GEN_679 ? registerTagMap_27_tagId : _GEN_706; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_708 = 5'h1c == _GEN_679 ? registerTagMap_28_tagId : _GEN_707; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_709 = 5'h1d == _GEN_679 ? registerTagMap_29_tagId : _GEN_708; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_710 = 5'h1e == _GEN_679 ? registerTagMap_30_tagId : _GEN_709; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_711 = 5'h1f == _GEN_679 ? registerTagMap_31_tagId : _GEN_710; // @[ReorderBuffer.scala 93:{17,17}]
  wire  _T_5 = index_2 == _GEN_711; // @[ReorderBuffer.scala 93:17]
  wire  _GEN_745 = 5'h1 == _GEN_679 ? 1'h0 : _GEN_547; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_746 = 5'h2 == _GEN_679 ? 1'h0 : _GEN_548; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_747 = 5'h3 == _GEN_679 ? 1'h0 : _GEN_549; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_748 = 5'h4 == _GEN_679 ? 1'h0 : _GEN_550; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_749 = 5'h5 == _GEN_679 ? 1'h0 : _GEN_551; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_750 = 5'h6 == _GEN_679 ? 1'h0 : _GEN_552; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_751 = 5'h7 == _GEN_679 ? 1'h0 : _GEN_553; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_752 = 5'h8 == _GEN_679 ? 1'h0 : _GEN_554; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_753 = 5'h9 == _GEN_679 ? 1'h0 : _GEN_555; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_754 = 5'ha == _GEN_679 ? 1'h0 : _GEN_556; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_755 = 5'hb == _GEN_679 ? 1'h0 : _GEN_557; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_756 = 5'hc == _GEN_679 ? 1'h0 : _GEN_558; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_757 = 5'hd == _GEN_679 ? 1'h0 : _GEN_559; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_758 = 5'he == _GEN_679 ? 1'h0 : _GEN_560; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_759 = 5'hf == _GEN_679 ? 1'h0 : _GEN_561; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_760 = 5'h10 == _GEN_679 ? 1'h0 : _GEN_562; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_761 = 5'h11 == _GEN_679 ? 1'h0 : _GEN_563; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_762 = 5'h12 == _GEN_679 ? 1'h0 : _GEN_564; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_763 = 5'h13 == _GEN_679 ? 1'h0 : _GEN_565; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_764 = 5'h14 == _GEN_679 ? 1'h0 : _GEN_566; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_765 = 5'h15 == _GEN_679 ? 1'h0 : _GEN_567; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_766 = 5'h16 == _GEN_679 ? 1'h0 : _GEN_568; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_767 = 5'h17 == _GEN_679 ? 1'h0 : _GEN_569; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_768 = 5'h18 == _GEN_679 ? 1'h0 : _GEN_570; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_769 = 5'h19 == _GEN_679 ? 1'h0 : _GEN_571; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_770 = 5'h1a == _GEN_679 ? 1'h0 : _GEN_572; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_771 = 5'h1b == _GEN_679 ? 1'h0 : _GEN_573; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_772 = 5'h1c == _GEN_679 ? 1'h0 : _GEN_574; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_773 = 5'h1d == _GEN_679 ? 1'h0 : _GEN_575; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_774 = 5'h1e == _GEN_679 ? 1'h0 : _GEN_576; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_775 = 5'h1f == _GEN_679 ? 1'h0 : _GEN_577; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_777 = _T_5 ? _GEN_745 : _GEN_547; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_778 = _T_5 ? _GEN_746 : _GEN_548; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_779 = _T_5 ? _GEN_747 : _GEN_549; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_780 = _T_5 ? _GEN_748 : _GEN_550; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_781 = _T_5 ? _GEN_749 : _GEN_551; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_782 = _T_5 ? _GEN_750 : _GEN_552; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_783 = _T_5 ? _GEN_751 : _GEN_553; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_784 = _T_5 ? _GEN_752 : _GEN_554; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_785 = _T_5 ? _GEN_753 : _GEN_555; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_786 = _T_5 ? _GEN_754 : _GEN_556; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_787 = _T_5 ? _GEN_755 : _GEN_557; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_788 = _T_5 ? _GEN_756 : _GEN_558; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_789 = _T_5 ? _GEN_757 : _GEN_559; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_790 = _T_5 ? _GEN_758 : _GEN_560; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_791 = _T_5 ? _GEN_759 : _GEN_561; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_792 = _T_5 ? _GEN_760 : _GEN_562; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_793 = _T_5 ? _GEN_761 : _GEN_563; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_794 = _T_5 ? _GEN_762 : _GEN_564; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_795 = _T_5 ? _GEN_763 : _GEN_565; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_796 = _T_5 ? _GEN_764 : _GEN_566; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_797 = _T_5 ? _GEN_765 : _GEN_567; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_798 = _T_5 ? _GEN_766 : _GEN_568; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_799 = _T_5 ? _GEN_767 : _GEN_569; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_800 = _T_5 ? _GEN_768 : _GEN_570; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_801 = _T_5 ? _GEN_769 : _GEN_571; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_802 = _T_5 ? _GEN_770 : _GEN_572; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_803 = _T_5 ? _GEN_771 : _GEN_573; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_804 = _T_5 ? _GEN_772 : _GEN_574; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_805 = _T_5 ? _GEN_773 : _GEN_575; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_806 = _T_5 ? _GEN_774 : _GEN_576; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_807 = _T_5 ? _GEN_775 : _GEN_577; // @[ReorderBuffer.scala 94:11]
  wire [63:0] _GEN_808 = _io_registerFile_2_valid_T ? _GEN_663 : 64'h0; // @[ReorderBuffer.scala 84:19 89:22 90:23]
  wire [4:0] _GEN_809 = _io_registerFile_2_valid_T ? _GEN_679 : 5'h0; // @[ReorderBuffer.scala 89:22 85:33 91:37]
  wire  _GEN_811 = _io_registerFile_2_valid_T ? _GEN_777 : _GEN_547; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_812 = _io_registerFile_2_valid_T ? _GEN_778 : _GEN_548; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_813 = _io_registerFile_2_valid_T ? _GEN_779 : _GEN_549; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_814 = _io_registerFile_2_valid_T ? _GEN_780 : _GEN_550; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_815 = _io_registerFile_2_valid_T ? _GEN_781 : _GEN_551; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_816 = _io_registerFile_2_valid_T ? _GEN_782 : _GEN_552; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_817 = _io_registerFile_2_valid_T ? _GEN_783 : _GEN_553; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_818 = _io_registerFile_2_valid_T ? _GEN_784 : _GEN_554; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_819 = _io_registerFile_2_valid_T ? _GEN_785 : _GEN_555; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_820 = _io_registerFile_2_valid_T ? _GEN_786 : _GEN_556; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_821 = _io_registerFile_2_valid_T ? _GEN_787 : _GEN_557; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_822 = _io_registerFile_2_valid_T ? _GEN_788 : _GEN_558; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_823 = _io_registerFile_2_valid_T ? _GEN_789 : _GEN_559; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_824 = _io_registerFile_2_valid_T ? _GEN_790 : _GEN_560; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_825 = _io_registerFile_2_valid_T ? _GEN_791 : _GEN_561; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_826 = _io_registerFile_2_valid_T ? _GEN_792 : _GEN_562; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_827 = _io_registerFile_2_valid_T ? _GEN_793 : _GEN_563; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_828 = _io_registerFile_2_valid_T ? _GEN_794 : _GEN_564; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_829 = _io_registerFile_2_valid_T ? _GEN_795 : _GEN_565; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_830 = _io_registerFile_2_valid_T ? _GEN_796 : _GEN_566; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_831 = _io_registerFile_2_valid_T ? _GEN_797 : _GEN_567; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_832 = _io_registerFile_2_valid_T ? _GEN_798 : _GEN_568; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_833 = _io_registerFile_2_valid_T ? _GEN_799 : _GEN_569; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_834 = _io_registerFile_2_valid_T ? _GEN_800 : _GEN_570; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_835 = _io_registerFile_2_valid_T ? _GEN_801 : _GEN_571; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_836 = _io_registerFile_2_valid_T ? _GEN_802 : _GEN_572; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_837 = _io_registerFile_2_valid_T ? _GEN_803 : _GEN_573; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_838 = _io_registerFile_2_valid_T ? _GEN_804 : _GEN_574; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_839 = _io_registerFile_2_valid_T ? _GEN_805 : _GEN_575; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_840 = _io_registerFile_2_valid_T ? _GEN_806 : _GEN_576; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_841 = _io_registerFile_2_valid_T ? _GEN_807 : _GEN_577; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_844 = _io_registerFile_2_valid_T ? _GEN_580 : 1'h1; // @[ReorderBuffer.scala 102:20 89:22]
  wire  _GEN_848 = canCommit_2 ? _GEN_811 : _GEN_547; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_849 = canCommit_2 ? _GEN_812 : _GEN_548; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_850 = canCommit_2 ? _GEN_813 : _GEN_549; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_851 = canCommit_2 ? _GEN_814 : _GEN_550; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_852 = canCommit_2 ? _GEN_815 : _GEN_551; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_853 = canCommit_2 ? _GEN_816 : _GEN_552; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_854 = canCommit_2 ? _GEN_817 : _GEN_553; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_855 = canCommit_2 ? _GEN_818 : _GEN_554; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_856 = canCommit_2 ? _GEN_819 : _GEN_555; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_857 = canCommit_2 ? _GEN_820 : _GEN_556; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_858 = canCommit_2 ? _GEN_821 : _GEN_557; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_859 = canCommit_2 ? _GEN_822 : _GEN_558; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_860 = canCommit_2 ? _GEN_823 : _GEN_559; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_861 = canCommit_2 ? _GEN_824 : _GEN_560; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_862 = canCommit_2 ? _GEN_825 : _GEN_561; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_863 = canCommit_2 ? _GEN_826 : _GEN_562; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_864 = canCommit_2 ? _GEN_827 : _GEN_563; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_865 = canCommit_2 ? _GEN_828 : _GEN_564; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_866 = canCommit_2 ? _GEN_829 : _GEN_565; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_867 = canCommit_2 ? _GEN_830 : _GEN_566; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_868 = canCommit_2 ? _GEN_831 : _GEN_567; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_869 = canCommit_2 ? _GEN_832 : _GEN_568; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_870 = canCommit_2 ? _GEN_833 : _GEN_569; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_871 = canCommit_2 ? _GEN_834 : _GEN_570; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_872 = canCommit_2 ? _GEN_835 : _GEN_571; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_873 = canCommit_2 ? _GEN_836 : _GEN_572; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_874 = canCommit_2 ? _GEN_837 : _GEN_573; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_875 = canCommit_2 ? _GEN_838 : _GEN_574; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_876 = canCommit_2 ? _GEN_839 : _GEN_575; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_877 = canCommit_2 ? _GEN_840 : _GEN_576; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_878 = canCommit_2 ? _GEN_841 : _GEN_577; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_881 = canCommit_2 ? _GEN_844 : _GEN_580; // @[ReorderBuffer.scala 88:21]
  wire [3:0] index_3 = tail + 4'h3; // @[ReorderBuffer.scala 77:22]
  wire  _GEN_902 = 4'h1 == index_3 ? buffer_1_valueReady : buffer_0_valueReady; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_903 = 4'h2 == index_3 ? buffer_2_valueReady : _GEN_902; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_904 = 4'h3 == index_3 ? buffer_3_valueReady : _GEN_903; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_905 = 4'h4 == index_3 ? buffer_4_valueReady : _GEN_904; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_906 = 4'h5 == index_3 ? buffer_5_valueReady : _GEN_905; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_907 = 4'h6 == index_3 ? buffer_6_valueReady : _GEN_906; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_908 = 4'h7 == index_3 ? buffer_7_valueReady : _GEN_907; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_909 = 4'h8 == index_3 ? buffer_8_valueReady : _GEN_908; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_910 = 4'h9 == index_3 ? buffer_9_valueReady : _GEN_909; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_911 = 4'ha == index_3 ? buffer_10_valueReady : _GEN_910; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_912 = 4'hb == index_3 ? buffer_11_valueReady : _GEN_911; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_913 = 4'hc == index_3 ? buffer_12_valueReady : _GEN_912; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_914 = 4'hd == index_3 ? buffer_13_valueReady : _GEN_913; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_915 = 4'he == index_3 ? buffer_14_valueReady : _GEN_914; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_916 = 4'hf == index_3 ? buffer_15_valueReady : _GEN_915; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_918 = 4'h1 == index_3 ? buffer_1_storeSign : buffer_0_storeSign; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_919 = 4'h2 == index_3 ? buffer_2_storeSign : _GEN_918; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_920 = 4'h3 == index_3 ? buffer_3_storeSign : _GEN_919; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_921 = 4'h4 == index_3 ? buffer_4_storeSign : _GEN_920; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_922 = 4'h5 == index_3 ? buffer_5_storeSign : _GEN_921; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_923 = 4'h6 == index_3 ? buffer_6_storeSign : _GEN_922; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_924 = 4'h7 == index_3 ? buffer_7_storeSign : _GEN_923; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_925 = 4'h8 == index_3 ? buffer_8_storeSign : _GEN_924; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_926 = 4'h9 == index_3 ? buffer_9_storeSign : _GEN_925; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_927 = 4'ha == index_3 ? buffer_10_storeSign : _GEN_926; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_928 = 4'hb == index_3 ? buffer_11_storeSign : _GEN_927; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_929 = 4'hc == index_3 ? buffer_12_storeSign : _GEN_928; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_930 = 4'hd == index_3 ? buffer_13_storeSign : _GEN_929; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_931 = 4'he == index_3 ? buffer_14_storeSign : _GEN_930; // @[ReorderBuffer.scala 79:{50,50}]
  wire  _GEN_932 = 4'hf == index_3 ? buffer_15_storeSign : _GEN_931; // @[ReorderBuffer.scala 79:{50,50}]
  wire  instructionOk_3 = _GEN_916 | _GEN_932; // @[ReorderBuffer.scala 79:50]
  wire  canCommit_3 = canCommit_2 & index_3 != head & instructionOk_3; // @[ReorderBuffer.scala 80:49]
  wire  _GEN_934 = 4'h1 == index_3 ? buffer_1_isError : buffer_0_isError; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_935 = 4'h2 == index_3 ? buffer_2_isError : _GEN_934; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_936 = 4'h3 == index_3 ? buffer_3_isError : _GEN_935; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_937 = 4'h4 == index_3 ? buffer_4_isError : _GEN_936; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_938 = 4'h5 == index_3 ? buffer_5_isError : _GEN_937; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_939 = 4'h6 == index_3 ? buffer_6_isError : _GEN_938; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_940 = 4'h7 == index_3 ? buffer_7_isError : _GEN_939; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_941 = 4'h8 == index_3 ? buffer_8_isError : _GEN_940; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_942 = 4'h9 == index_3 ? buffer_9_isError : _GEN_941; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_943 = 4'ha == index_3 ? buffer_10_isError : _GEN_942; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_944 = 4'hb == index_3 ? buffer_11_isError : _GEN_943; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_945 = 4'hc == index_3 ? buffer_12_isError : _GEN_944; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_946 = 4'hd == index_3 ? buffer_13_isError : _GEN_945; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_947 = 4'he == index_3 ? buffer_14_isError : _GEN_946; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _GEN_948 = 4'hf == index_3 ? buffer_15_isError : _GEN_947; // @[ReorderBuffer.scala 83:{30,30}]
  wire  _io_registerFile_3_valid_T = ~_GEN_948; // @[ReorderBuffer.scala 83:30]
  wire [63:0] _GEN_950 = 4'h1 == index_3 ? buffer_1_value : buffer_0_value; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_951 = 4'h2 == index_3 ? buffer_2_value : _GEN_950; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_952 = 4'h3 == index_3 ? buffer_3_value : _GEN_951; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_953 = 4'h4 == index_3 ? buffer_4_value : _GEN_952; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_954 = 4'h5 == index_3 ? buffer_5_value : _GEN_953; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_955 = 4'h6 == index_3 ? buffer_6_value : _GEN_954; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_956 = 4'h7 == index_3 ? buffer_7_value : _GEN_955; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_957 = 4'h8 == index_3 ? buffer_8_value : _GEN_956; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_958 = 4'h9 == index_3 ? buffer_9_value : _GEN_957; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_959 = 4'ha == index_3 ? buffer_10_value : _GEN_958; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_960 = 4'hb == index_3 ? buffer_11_value : _GEN_959; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_961 = 4'hc == index_3 ? buffer_12_value : _GEN_960; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_962 = 4'hd == index_3 ? buffer_13_value : _GEN_961; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_963 = 4'he == index_3 ? buffer_14_value : _GEN_962; // @[ReorderBuffer.scala 90:{23,23}]
  wire [63:0] _GEN_964 = 4'hf == index_3 ? buffer_15_value : _GEN_963; // @[ReorderBuffer.scala 90:{23,23}]
  wire [4:0] _GEN_966 = 4'h1 == index_3 ? buffer_1_destinationRegister : buffer_0_destinationRegister; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_967 = 4'h2 == index_3 ? buffer_2_destinationRegister : _GEN_966; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_968 = 4'h3 == index_3 ? buffer_3_destinationRegister : _GEN_967; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_969 = 4'h4 == index_3 ? buffer_4_destinationRegister : _GEN_968; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_970 = 4'h5 == index_3 ? buffer_5_destinationRegister : _GEN_969; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_971 = 4'h6 == index_3 ? buffer_6_destinationRegister : _GEN_970; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_972 = 4'h7 == index_3 ? buffer_7_destinationRegister : _GEN_971; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_973 = 4'h8 == index_3 ? buffer_8_destinationRegister : _GEN_972; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_974 = 4'h9 == index_3 ? buffer_9_destinationRegister : _GEN_973; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_975 = 4'ha == index_3 ? buffer_10_destinationRegister : _GEN_974; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_976 = 4'hb == index_3 ? buffer_11_destinationRegister : _GEN_975; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_977 = 4'hc == index_3 ? buffer_12_destinationRegister : _GEN_976; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_978 = 4'hd == index_3 ? buffer_13_destinationRegister : _GEN_977; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_979 = 4'he == index_3 ? buffer_14_destinationRegister : _GEN_978; // @[ReorderBuffer.scala 91:{37,37}]
  wire [4:0] _GEN_980 = 4'hf == index_3 ? buffer_15_destinationRegister : _GEN_979; // @[ReorderBuffer.scala 91:{37,37}]
  wire [3:0] _GEN_982 = 5'h1 == _GEN_980 ? registerTagMap_1_tagId : 4'h0; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_983 = 5'h2 == _GEN_980 ? registerTagMap_2_tagId : _GEN_982; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_984 = 5'h3 == _GEN_980 ? registerTagMap_3_tagId : _GEN_983; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_985 = 5'h4 == _GEN_980 ? registerTagMap_4_tagId : _GEN_984; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_986 = 5'h5 == _GEN_980 ? registerTagMap_5_tagId : _GEN_985; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_987 = 5'h6 == _GEN_980 ? registerTagMap_6_tagId : _GEN_986; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_988 = 5'h7 == _GEN_980 ? registerTagMap_7_tagId : _GEN_987; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_989 = 5'h8 == _GEN_980 ? registerTagMap_8_tagId : _GEN_988; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_990 = 5'h9 == _GEN_980 ? registerTagMap_9_tagId : _GEN_989; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_991 = 5'ha == _GEN_980 ? registerTagMap_10_tagId : _GEN_990; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_992 = 5'hb == _GEN_980 ? registerTagMap_11_tagId : _GEN_991; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_993 = 5'hc == _GEN_980 ? registerTagMap_12_tagId : _GEN_992; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_994 = 5'hd == _GEN_980 ? registerTagMap_13_tagId : _GEN_993; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_995 = 5'he == _GEN_980 ? registerTagMap_14_tagId : _GEN_994; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_996 = 5'hf == _GEN_980 ? registerTagMap_15_tagId : _GEN_995; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_997 = 5'h10 == _GEN_980 ? registerTagMap_16_tagId : _GEN_996; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_998 = 5'h11 == _GEN_980 ? registerTagMap_17_tagId : _GEN_997; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_999 = 5'h12 == _GEN_980 ? registerTagMap_18_tagId : _GEN_998; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_1000 = 5'h13 == _GEN_980 ? registerTagMap_19_tagId : _GEN_999; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_1001 = 5'h14 == _GEN_980 ? registerTagMap_20_tagId : _GEN_1000; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_1002 = 5'h15 == _GEN_980 ? registerTagMap_21_tagId : _GEN_1001; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_1003 = 5'h16 == _GEN_980 ? registerTagMap_22_tagId : _GEN_1002; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_1004 = 5'h17 == _GEN_980 ? registerTagMap_23_tagId : _GEN_1003; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_1005 = 5'h18 == _GEN_980 ? registerTagMap_24_tagId : _GEN_1004; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_1006 = 5'h19 == _GEN_980 ? registerTagMap_25_tagId : _GEN_1005; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_1007 = 5'h1a == _GEN_980 ? registerTagMap_26_tagId : _GEN_1006; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_1008 = 5'h1b == _GEN_980 ? registerTagMap_27_tagId : _GEN_1007; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_1009 = 5'h1c == _GEN_980 ? registerTagMap_28_tagId : _GEN_1008; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_1010 = 5'h1d == _GEN_980 ? registerTagMap_29_tagId : _GEN_1009; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_1011 = 5'h1e == _GEN_980 ? registerTagMap_30_tagId : _GEN_1010; // @[ReorderBuffer.scala 93:{17,17}]
  wire [3:0] _GEN_1012 = 5'h1f == _GEN_980 ? registerTagMap_31_tagId : _GEN_1011; // @[ReorderBuffer.scala 93:{17,17}]
  wire  _T_7 = index_3 == _GEN_1012; // @[ReorderBuffer.scala 93:17]
  wire  _GEN_1046 = 5'h1 == _GEN_980 ? 1'h0 : _GEN_848; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_1047 = 5'h2 == _GEN_980 ? 1'h0 : _GEN_849; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_1048 = 5'h3 == _GEN_980 ? 1'h0 : _GEN_850; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_1049 = 5'h4 == _GEN_980 ? 1'h0 : _GEN_851; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_1050 = 5'h5 == _GEN_980 ? 1'h0 : _GEN_852; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_1051 = 5'h6 == _GEN_980 ? 1'h0 : _GEN_853; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_1052 = 5'h7 == _GEN_980 ? 1'h0 : _GEN_854; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_1053 = 5'h8 == _GEN_980 ? 1'h0 : _GEN_855; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_1054 = 5'h9 == _GEN_980 ? 1'h0 : _GEN_856; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_1055 = 5'ha == _GEN_980 ? 1'h0 : _GEN_857; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_1056 = 5'hb == _GEN_980 ? 1'h0 : _GEN_858; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_1057 = 5'hc == _GEN_980 ? 1'h0 : _GEN_859; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_1058 = 5'hd == _GEN_980 ? 1'h0 : _GEN_860; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_1059 = 5'he == _GEN_980 ? 1'h0 : _GEN_861; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_1060 = 5'hf == _GEN_980 ? 1'h0 : _GEN_862; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_1061 = 5'h10 == _GEN_980 ? 1'h0 : _GEN_863; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_1062 = 5'h11 == _GEN_980 ? 1'h0 : _GEN_864; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_1063 = 5'h12 == _GEN_980 ? 1'h0 : _GEN_865; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_1064 = 5'h13 == _GEN_980 ? 1'h0 : _GEN_866; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_1065 = 5'h14 == _GEN_980 ? 1'h0 : _GEN_867; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_1066 = 5'h15 == _GEN_980 ? 1'h0 : _GEN_868; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_1067 = 5'h16 == _GEN_980 ? 1'h0 : _GEN_869; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_1068 = 5'h17 == _GEN_980 ? 1'h0 : _GEN_870; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_1069 = 5'h18 == _GEN_980 ? 1'h0 : _GEN_871; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_1070 = 5'h19 == _GEN_980 ? 1'h0 : _GEN_872; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_1071 = 5'h1a == _GEN_980 ? 1'h0 : _GEN_873; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_1072 = 5'h1b == _GEN_980 ? 1'h0 : _GEN_874; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_1073 = 5'h1c == _GEN_980 ? 1'h0 : _GEN_875; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_1074 = 5'h1d == _GEN_980 ? 1'h0 : _GEN_876; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_1075 = 5'h1e == _GEN_980 ? 1'h0 : _GEN_877; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_1076 = 5'h1f == _GEN_980 ? 1'h0 : _GEN_878; // @[ReorderBuffer.scala 97:{13,13}]
  wire  _GEN_1078 = _T_7 ? _GEN_1046 : _GEN_848; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_1079 = _T_7 ? _GEN_1047 : _GEN_849; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_1080 = _T_7 ? _GEN_1048 : _GEN_850; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_1081 = _T_7 ? _GEN_1049 : _GEN_851; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_1082 = _T_7 ? _GEN_1050 : _GEN_852; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_1083 = _T_7 ? _GEN_1051 : _GEN_853; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_1084 = _T_7 ? _GEN_1052 : _GEN_854; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_1085 = _T_7 ? _GEN_1053 : _GEN_855; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_1086 = _T_7 ? _GEN_1054 : _GEN_856; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_1087 = _T_7 ? _GEN_1055 : _GEN_857; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_1088 = _T_7 ? _GEN_1056 : _GEN_858; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_1089 = _T_7 ? _GEN_1057 : _GEN_859; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_1090 = _T_7 ? _GEN_1058 : _GEN_860; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_1091 = _T_7 ? _GEN_1059 : _GEN_861; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_1092 = _T_7 ? _GEN_1060 : _GEN_862; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_1093 = _T_7 ? _GEN_1061 : _GEN_863; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_1094 = _T_7 ? _GEN_1062 : _GEN_864; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_1095 = _T_7 ? _GEN_1063 : _GEN_865; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_1096 = _T_7 ? _GEN_1064 : _GEN_866; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_1097 = _T_7 ? _GEN_1065 : _GEN_867; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_1098 = _T_7 ? _GEN_1066 : _GEN_868; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_1099 = _T_7 ? _GEN_1067 : _GEN_869; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_1100 = _T_7 ? _GEN_1068 : _GEN_870; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_1101 = _T_7 ? _GEN_1069 : _GEN_871; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_1102 = _T_7 ? _GEN_1070 : _GEN_872; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_1103 = _T_7 ? _GEN_1071 : _GEN_873; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_1104 = _T_7 ? _GEN_1072 : _GEN_874; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_1105 = _T_7 ? _GEN_1073 : _GEN_875; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_1106 = _T_7 ? _GEN_1074 : _GEN_876; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_1107 = _T_7 ? _GEN_1075 : _GEN_877; // @[ReorderBuffer.scala 94:11]
  wire  _GEN_1108 = _T_7 ? _GEN_1076 : _GEN_878; // @[ReorderBuffer.scala 94:11]
  wire [63:0] _GEN_1109 = _io_registerFile_3_valid_T ? _GEN_964 : 64'h0; // @[ReorderBuffer.scala 84:19 89:22 90:23]
  wire [4:0] _GEN_1110 = _io_registerFile_3_valid_T ? _GEN_980 : 5'h0; // @[ReorderBuffer.scala 89:22 85:33 91:37]
  wire  _GEN_1112 = _io_registerFile_3_valid_T ? _GEN_1078 : _GEN_848; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_1113 = _io_registerFile_3_valid_T ? _GEN_1079 : _GEN_849; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_1114 = _io_registerFile_3_valid_T ? _GEN_1080 : _GEN_850; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_1115 = _io_registerFile_3_valid_T ? _GEN_1081 : _GEN_851; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_1116 = _io_registerFile_3_valid_T ? _GEN_1082 : _GEN_852; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_1117 = _io_registerFile_3_valid_T ? _GEN_1083 : _GEN_853; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_1118 = _io_registerFile_3_valid_T ? _GEN_1084 : _GEN_854; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_1119 = _io_registerFile_3_valid_T ? _GEN_1085 : _GEN_855; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_1120 = _io_registerFile_3_valid_T ? _GEN_1086 : _GEN_856; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_1121 = _io_registerFile_3_valid_T ? _GEN_1087 : _GEN_857; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_1122 = _io_registerFile_3_valid_T ? _GEN_1088 : _GEN_858; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_1123 = _io_registerFile_3_valid_T ? _GEN_1089 : _GEN_859; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_1124 = _io_registerFile_3_valid_T ? _GEN_1090 : _GEN_860; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_1125 = _io_registerFile_3_valid_T ? _GEN_1091 : _GEN_861; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_1126 = _io_registerFile_3_valid_T ? _GEN_1092 : _GEN_862; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_1127 = _io_registerFile_3_valid_T ? _GEN_1093 : _GEN_863; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_1128 = _io_registerFile_3_valid_T ? _GEN_1094 : _GEN_864; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_1129 = _io_registerFile_3_valid_T ? _GEN_1095 : _GEN_865; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_1130 = _io_registerFile_3_valid_T ? _GEN_1096 : _GEN_866; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_1131 = _io_registerFile_3_valid_T ? _GEN_1097 : _GEN_867; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_1132 = _io_registerFile_3_valid_T ? _GEN_1098 : _GEN_868; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_1133 = _io_registerFile_3_valid_T ? _GEN_1099 : _GEN_869; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_1134 = _io_registerFile_3_valid_T ? _GEN_1100 : _GEN_870; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_1135 = _io_registerFile_3_valid_T ? _GEN_1101 : _GEN_871; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_1136 = _io_registerFile_3_valid_T ? _GEN_1102 : _GEN_872; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_1137 = _io_registerFile_3_valid_T ? _GEN_1103 : _GEN_873; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_1138 = _io_registerFile_3_valid_T ? _GEN_1104 : _GEN_874; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_1139 = _io_registerFile_3_valid_T ? _GEN_1105 : _GEN_875; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_1140 = _io_registerFile_3_valid_T ? _GEN_1106 : _GEN_876; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_1141 = _io_registerFile_3_valid_T ? _GEN_1107 : _GEN_877; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_1142 = _io_registerFile_3_valid_T ? _GEN_1108 : _GEN_878; // @[ReorderBuffer.scala 89:22]
  wire  _GEN_1145 = _io_registerFile_3_valid_T ? _GEN_881 : 1'h1; // @[ReorderBuffer.scala 102:20 89:22]
  wire  _GEN_1149 = canCommit_3 ? _GEN_1112 : _GEN_848; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_1150 = canCommit_3 ? _GEN_1113 : _GEN_849; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_1151 = canCommit_3 ? _GEN_1114 : _GEN_850; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_1152 = canCommit_3 ? _GEN_1115 : _GEN_851; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_1153 = canCommit_3 ? _GEN_1116 : _GEN_852; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_1154 = canCommit_3 ? _GEN_1117 : _GEN_853; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_1155 = canCommit_3 ? _GEN_1118 : _GEN_854; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_1156 = canCommit_3 ? _GEN_1119 : _GEN_855; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_1157 = canCommit_3 ? _GEN_1120 : _GEN_856; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_1158 = canCommit_3 ? _GEN_1121 : _GEN_857; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_1159 = canCommit_3 ? _GEN_1122 : _GEN_858; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_1160 = canCommit_3 ? _GEN_1123 : _GEN_859; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_1161 = canCommit_3 ? _GEN_1124 : _GEN_860; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_1162 = canCommit_3 ? _GEN_1125 : _GEN_861; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_1163 = canCommit_3 ? _GEN_1126 : _GEN_862; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_1164 = canCommit_3 ? _GEN_1127 : _GEN_863; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_1165 = canCommit_3 ? _GEN_1128 : _GEN_864; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_1166 = canCommit_3 ? _GEN_1129 : _GEN_865; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_1167 = canCommit_3 ? _GEN_1130 : _GEN_866; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_1168 = canCommit_3 ? _GEN_1131 : _GEN_867; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_1169 = canCommit_3 ? _GEN_1132 : _GEN_868; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_1170 = canCommit_3 ? _GEN_1133 : _GEN_869; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_1171 = canCommit_3 ? _GEN_1134 : _GEN_870; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_1172 = canCommit_3 ? _GEN_1135 : _GEN_871; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_1173 = canCommit_3 ? _GEN_1136 : _GEN_872; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_1174 = canCommit_3 ? _GEN_1137 : _GEN_873; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_1175 = canCommit_3 ? _GEN_1138 : _GEN_874; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_1176 = canCommit_3 ? _GEN_1139 : _GEN_875; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_1177 = canCommit_3 ? _GEN_1140 : _GEN_876; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_1178 = canCommit_3 ? _GEN_1141 : _GEN_877; // @[ReorderBuffer.scala 88:21]
  wire  _GEN_1179 = canCommit_3 ? _GEN_1142 : _GEN_878; // @[ReorderBuffer.scala 88:21]
  wire  _tailDelta_T = ~io_registerFile_0_valid; // @[ReorderBuffer.scala 120:7]
  wire  _tailDelta_T_1 = ~io_registerFile_1_valid; // @[ReorderBuffer.scala 120:7]
  wire  _tailDelta_T_2 = ~io_registerFile_2_valid; // @[ReorderBuffer.scala 120:7]
  wire  _tailDelta_T_3 = ~io_registerFile_3_valid; // @[ReorderBuffer.scala 120:7]
  wire [2:0] _tailDelta_T_4 = _tailDelta_T_3 ? 3'h3 : 3'h4; // @[Mux.scala 101:16]
  wire [2:0] _tailDelta_T_5 = _tailDelta_T_2 ? 3'h2 : _tailDelta_T_4; // @[Mux.scala 101:16]
  wire [2:0] _tailDelta_T_6 = _tailDelta_T_1 ? 3'h1 : _tailDelta_T_5; // @[Mux.scala 101:16]
  wire [2:0] tailDelta = _tailDelta_T ? 3'h0 : _tailDelta_T_6; // @[Mux.scala 101:16]
  wire [3:0] _io_decoders_0_ready_T_1 = head + 4'h1; // @[ReorderBuffer.scala 129:48]
  wire  _T_8 = io_decoders_0_valid & io_decoders_0_ready; // @[ReorderBuffer.scala 130:24]
  wire  _GEN_1218 = 4'h0 == head ? 1'h0 : buffer_0_valueReady; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire  _GEN_1219 = 4'h1 == head ? 1'h0 : buffer_1_valueReady; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire  _GEN_1220 = 4'h2 == head ? 1'h0 : buffer_2_valueReady; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire  _GEN_1221 = 4'h3 == head ? 1'h0 : buffer_3_valueReady; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire  _GEN_1222 = 4'h4 == head ? 1'h0 : buffer_4_valueReady; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire  _GEN_1223 = 4'h5 == head ? 1'h0 : buffer_5_valueReady; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire  _GEN_1224 = 4'h6 == head ? 1'h0 : buffer_6_valueReady; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire  _GEN_1225 = 4'h7 == head ? 1'h0 : buffer_7_valueReady; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire  _GEN_1226 = 4'h8 == head ? 1'h0 : buffer_8_valueReady; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire  _GEN_1227 = 4'h9 == head ? 1'h0 : buffer_9_valueReady; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire  _GEN_1228 = 4'ha == head ? 1'h0 : buffer_10_valueReady; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire  _GEN_1229 = 4'hb == head ? 1'h0 : buffer_11_valueReady; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire  _GEN_1230 = 4'hc == head ? 1'h0 : buffer_12_valueReady; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire  _GEN_1231 = 4'hd == head ? 1'h0 : buffer_13_valueReady; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire  _GEN_1232 = 4'he == head ? 1'h0 : buffer_14_valueReady; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire  _GEN_1233 = 4'hf == head ? 1'h0 : buffer_15_valueReady; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire [63:0] _GEN_1234 = 4'h0 == head ? 64'h0 : buffer_0_value; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire [63:0] _GEN_1235 = 4'h1 == head ? 64'h0 : buffer_1_value; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire [63:0] _GEN_1236 = 4'h2 == head ? 64'h0 : buffer_2_value; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire [63:0] _GEN_1237 = 4'h3 == head ? 64'h0 : buffer_3_value; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire [63:0] _GEN_1238 = 4'h4 == head ? 64'h0 : buffer_4_value; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire [63:0] _GEN_1239 = 4'h5 == head ? 64'h0 : buffer_5_value; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire [63:0] _GEN_1240 = 4'h6 == head ? 64'h0 : buffer_6_value; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire [63:0] _GEN_1241 = 4'h7 == head ? 64'h0 : buffer_7_value; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire [63:0] _GEN_1242 = 4'h8 == head ? 64'h0 : buffer_8_value; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire [63:0] _GEN_1243 = 4'h9 == head ? 64'h0 : buffer_9_value; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire [63:0] _GEN_1244 = 4'ha == head ? 64'h0 : buffer_10_value; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire [63:0] _GEN_1245 = 4'hb == head ? 64'h0 : buffer_11_value; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire [63:0] _GEN_1246 = 4'hc == head ? 64'h0 : buffer_12_value; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire [63:0] _GEN_1247 = 4'hd == head ? 64'h0 : buffer_13_value; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire [63:0] _GEN_1248 = 4'he == head ? 64'h0 : buffer_14_value; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire [63:0] _GEN_1249 = 4'hf == head ? 64'h0 : buffer_15_value; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire  _GEN_1282 = 4'h0 == head ? 1'h0 : buffer_0_isError; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire  _GEN_1283 = 4'h1 == head ? 1'h0 : buffer_1_isError; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire  _GEN_1284 = 4'h2 == head ? 1'h0 : buffer_2_isError; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire  _GEN_1285 = 4'h3 == head ? 1'h0 : buffer_3_isError; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire  _GEN_1286 = 4'h4 == head ? 1'h0 : buffer_4_isError; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire  _GEN_1287 = 4'h5 == head ? 1'h0 : buffer_5_isError; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire  _GEN_1288 = 4'h6 == head ? 1'h0 : buffer_6_isError; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire  _GEN_1289 = 4'h7 == head ? 1'h0 : buffer_7_isError; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire  _GEN_1290 = 4'h8 == head ? 1'h0 : buffer_8_isError; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire  _GEN_1291 = 4'h9 == head ? 1'h0 : buffer_9_isError; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire  _GEN_1292 = 4'ha == head ? 1'h0 : buffer_10_isError; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire  _GEN_1293 = 4'hb == head ? 1'h0 : buffer_11_isError; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire  _GEN_1294 = 4'hc == head ? 1'h0 : buffer_12_isError; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire  _GEN_1295 = 4'hd == head ? 1'h0 : buffer_13_isError; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire  _GEN_1296 = 4'he == head ? 1'h0 : buffer_14_isError; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire  _GEN_1297 = 4'hf == head ? 1'h0 : buffer_15_isError; // @[ReorderBuffer.scala 133:{27,27} 55:23]
  wire  _GEN_1314 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1218 : buffer_0_valueReady; // @[ReorderBuffer.scala 130:42 55:23]
  wire  _GEN_1315 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1219 : buffer_1_valueReady; // @[ReorderBuffer.scala 130:42 55:23]
  wire  _GEN_1316 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1220 : buffer_2_valueReady; // @[ReorderBuffer.scala 130:42 55:23]
  wire  _GEN_1317 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1221 : buffer_3_valueReady; // @[ReorderBuffer.scala 130:42 55:23]
  wire  _GEN_1318 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1222 : buffer_4_valueReady; // @[ReorderBuffer.scala 130:42 55:23]
  wire  _GEN_1319 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1223 : buffer_5_valueReady; // @[ReorderBuffer.scala 130:42 55:23]
  wire  _GEN_1320 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1224 : buffer_6_valueReady; // @[ReorderBuffer.scala 130:42 55:23]
  wire  _GEN_1321 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1225 : buffer_7_valueReady; // @[ReorderBuffer.scala 130:42 55:23]
  wire  _GEN_1322 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1226 : buffer_8_valueReady; // @[ReorderBuffer.scala 130:42 55:23]
  wire  _GEN_1323 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1227 : buffer_9_valueReady; // @[ReorderBuffer.scala 130:42 55:23]
  wire  _GEN_1324 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1228 : buffer_10_valueReady; // @[ReorderBuffer.scala 130:42 55:23]
  wire  _GEN_1325 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1229 : buffer_11_valueReady; // @[ReorderBuffer.scala 130:42 55:23]
  wire  _GEN_1326 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1230 : buffer_12_valueReady; // @[ReorderBuffer.scala 130:42 55:23]
  wire  _GEN_1327 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1231 : buffer_13_valueReady; // @[ReorderBuffer.scala 130:42 55:23]
  wire  _GEN_1328 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1232 : buffer_14_valueReady; // @[ReorderBuffer.scala 130:42 55:23]
  wire  _GEN_1329 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1233 : buffer_15_valueReady; // @[ReorderBuffer.scala 130:42 55:23]
  wire [63:0] _GEN_1330 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1234 : buffer_0_value; // @[ReorderBuffer.scala 130:42 55:23]
  wire [63:0] _GEN_1331 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1235 : buffer_1_value; // @[ReorderBuffer.scala 130:42 55:23]
  wire [63:0] _GEN_1332 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1236 : buffer_2_value; // @[ReorderBuffer.scala 130:42 55:23]
  wire [63:0] _GEN_1333 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1237 : buffer_3_value; // @[ReorderBuffer.scala 130:42 55:23]
  wire [63:0] _GEN_1334 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1238 : buffer_4_value; // @[ReorderBuffer.scala 130:42 55:23]
  wire [63:0] _GEN_1335 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1239 : buffer_5_value; // @[ReorderBuffer.scala 130:42 55:23]
  wire [63:0] _GEN_1336 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1240 : buffer_6_value; // @[ReorderBuffer.scala 130:42 55:23]
  wire [63:0] _GEN_1337 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1241 : buffer_7_value; // @[ReorderBuffer.scala 130:42 55:23]
  wire [63:0] _GEN_1338 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1242 : buffer_8_value; // @[ReorderBuffer.scala 130:42 55:23]
  wire [63:0] _GEN_1339 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1243 : buffer_9_value; // @[ReorderBuffer.scala 130:42 55:23]
  wire [63:0] _GEN_1340 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1244 : buffer_10_value; // @[ReorderBuffer.scala 130:42 55:23]
  wire [63:0] _GEN_1341 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1245 : buffer_11_value; // @[ReorderBuffer.scala 130:42 55:23]
  wire [63:0] _GEN_1342 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1246 : buffer_12_value; // @[ReorderBuffer.scala 130:42 55:23]
  wire [63:0] _GEN_1343 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1247 : buffer_13_value; // @[ReorderBuffer.scala 130:42 55:23]
  wire [63:0] _GEN_1344 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1248 : buffer_14_value; // @[ReorderBuffer.scala 130:42 55:23]
  wire [63:0] _GEN_1345 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1249 : buffer_15_value; // @[ReorderBuffer.scala 130:42 55:23]
  wire  _GEN_1378 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1282 : buffer_0_isError; // @[ReorderBuffer.scala 130:42 55:23]
  wire  _GEN_1379 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1283 : buffer_1_isError; // @[ReorderBuffer.scala 130:42 55:23]
  wire  _GEN_1380 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1284 : buffer_2_isError; // @[ReorderBuffer.scala 130:42 55:23]
  wire  _GEN_1381 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1285 : buffer_3_isError; // @[ReorderBuffer.scala 130:42 55:23]
  wire  _GEN_1382 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1286 : buffer_4_isError; // @[ReorderBuffer.scala 130:42 55:23]
  wire  _GEN_1383 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1287 : buffer_5_isError; // @[ReorderBuffer.scala 130:42 55:23]
  wire  _GEN_1384 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1288 : buffer_6_isError; // @[ReorderBuffer.scala 130:42 55:23]
  wire  _GEN_1385 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1289 : buffer_7_isError; // @[ReorderBuffer.scala 130:42 55:23]
  wire  _GEN_1386 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1290 : buffer_8_isError; // @[ReorderBuffer.scala 130:42 55:23]
  wire  _GEN_1387 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1291 : buffer_9_isError; // @[ReorderBuffer.scala 130:42 55:23]
  wire  _GEN_1388 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1292 : buffer_10_isError; // @[ReorderBuffer.scala 130:42 55:23]
  wire  _GEN_1389 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1293 : buffer_11_isError; // @[ReorderBuffer.scala 130:42 55:23]
  wire  _GEN_1390 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1294 : buffer_12_isError; // @[ReorderBuffer.scala 130:42 55:23]
  wire  _GEN_1391 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1295 : buffer_13_isError; // @[ReorderBuffer.scala 130:42 55:23]
  wire  _GEN_1392 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1296 : buffer_14_isError; // @[ReorderBuffer.scala 130:42 55:23]
  wire  _GEN_1393 = io_decoders_0_valid & io_decoders_0_ready ? _GEN_1297 : buffer_15_isError; // @[ReorderBuffer.scala 130:42 55:23]
  wire  _GEN_1395 = 5'h1 == io_decoders_0_destination_destinationRegister | _GEN_1149; // @[ReorderBuffer.scala 146:{69,69}]
  wire  _GEN_1396 = 5'h2 == io_decoders_0_destination_destinationRegister | _GEN_1150; // @[ReorderBuffer.scala 146:{69,69}]
  wire  _GEN_1397 = 5'h3 == io_decoders_0_destination_destinationRegister | _GEN_1151; // @[ReorderBuffer.scala 146:{69,69}]
  wire  _GEN_1398 = 5'h4 == io_decoders_0_destination_destinationRegister | _GEN_1152; // @[ReorderBuffer.scala 146:{69,69}]
  wire  _GEN_1399 = 5'h5 == io_decoders_0_destination_destinationRegister | _GEN_1153; // @[ReorderBuffer.scala 146:{69,69}]
  wire  _GEN_1400 = 5'h6 == io_decoders_0_destination_destinationRegister | _GEN_1154; // @[ReorderBuffer.scala 146:{69,69}]
  wire  _GEN_1401 = 5'h7 == io_decoders_0_destination_destinationRegister | _GEN_1155; // @[ReorderBuffer.scala 146:{69,69}]
  wire  _GEN_1402 = 5'h8 == io_decoders_0_destination_destinationRegister | _GEN_1156; // @[ReorderBuffer.scala 146:{69,69}]
  wire  _GEN_1403 = 5'h9 == io_decoders_0_destination_destinationRegister | _GEN_1157; // @[ReorderBuffer.scala 146:{69,69}]
  wire  _GEN_1404 = 5'ha == io_decoders_0_destination_destinationRegister | _GEN_1158; // @[ReorderBuffer.scala 146:{69,69}]
  wire  _GEN_1405 = 5'hb == io_decoders_0_destination_destinationRegister | _GEN_1159; // @[ReorderBuffer.scala 146:{69,69}]
  wire  _GEN_1406 = 5'hc == io_decoders_0_destination_destinationRegister | _GEN_1160; // @[ReorderBuffer.scala 146:{69,69}]
  wire  _GEN_1407 = 5'hd == io_decoders_0_destination_destinationRegister | _GEN_1161; // @[ReorderBuffer.scala 146:{69,69}]
  wire  _GEN_1408 = 5'he == io_decoders_0_destination_destinationRegister | _GEN_1162; // @[ReorderBuffer.scala 146:{69,69}]
  wire  _GEN_1409 = 5'hf == io_decoders_0_destination_destinationRegister | _GEN_1163; // @[ReorderBuffer.scala 146:{69,69}]
  wire  _GEN_1410 = 5'h10 == io_decoders_0_destination_destinationRegister | _GEN_1164; // @[ReorderBuffer.scala 146:{69,69}]
  wire  _GEN_1411 = 5'h11 == io_decoders_0_destination_destinationRegister | _GEN_1165; // @[ReorderBuffer.scala 146:{69,69}]
  wire  _GEN_1412 = 5'h12 == io_decoders_0_destination_destinationRegister | _GEN_1166; // @[ReorderBuffer.scala 146:{69,69}]
  wire  _GEN_1413 = 5'h13 == io_decoders_0_destination_destinationRegister | _GEN_1167; // @[ReorderBuffer.scala 146:{69,69}]
  wire  _GEN_1414 = 5'h14 == io_decoders_0_destination_destinationRegister | _GEN_1168; // @[ReorderBuffer.scala 146:{69,69}]
  wire  _GEN_1415 = 5'h15 == io_decoders_0_destination_destinationRegister | _GEN_1169; // @[ReorderBuffer.scala 146:{69,69}]
  wire  _GEN_1416 = 5'h16 == io_decoders_0_destination_destinationRegister | _GEN_1170; // @[ReorderBuffer.scala 146:{69,69}]
  wire  _GEN_1417 = 5'h17 == io_decoders_0_destination_destinationRegister | _GEN_1171; // @[ReorderBuffer.scala 146:{69,69}]
  wire  _GEN_1418 = 5'h18 == io_decoders_0_destination_destinationRegister | _GEN_1172; // @[ReorderBuffer.scala 146:{69,69}]
  wire  _GEN_1419 = 5'h19 == io_decoders_0_destination_destinationRegister | _GEN_1173; // @[ReorderBuffer.scala 146:{69,69}]
  wire  _GEN_1420 = 5'h1a == io_decoders_0_destination_destinationRegister | _GEN_1174; // @[ReorderBuffer.scala 146:{69,69}]
  wire  _GEN_1421 = 5'h1b == io_decoders_0_destination_destinationRegister | _GEN_1175; // @[ReorderBuffer.scala 146:{69,69}]
  wire  _GEN_1422 = 5'h1c == io_decoders_0_destination_destinationRegister | _GEN_1176; // @[ReorderBuffer.scala 146:{69,69}]
  wire  _GEN_1423 = 5'h1d == io_decoders_0_destination_destinationRegister | _GEN_1177; // @[ReorderBuffer.scala 146:{69,69}]
  wire  _GEN_1424 = 5'h1e == io_decoders_0_destination_destinationRegister | _GEN_1178; // @[ReorderBuffer.scala 146:{69,69}]
  wire  _GEN_1425 = 5'h1f == io_decoders_0_destination_destinationRegister | _GEN_1179; // @[ReorderBuffer.scala 146:{69,69}]
  wire  _GEN_1524 = 5'h2 == io_decoders_0_source1_sourceRegister ? registerTagMap_2_valid : 5'h1 ==
    io_decoders_0_source1_sourceRegister & registerTagMap_1_valid; // @[ReorderBuffer.scala 155:{41,41}]
  wire  _GEN_1525 = 5'h3 == io_decoders_0_source1_sourceRegister ? registerTagMap_3_valid : _GEN_1524; // @[ReorderBuffer.scala 155:{41,41}]
  wire  _GEN_1526 = 5'h4 == io_decoders_0_source1_sourceRegister ? registerTagMap_4_valid : _GEN_1525; // @[ReorderBuffer.scala 155:{41,41}]
  wire  _GEN_1527 = 5'h5 == io_decoders_0_source1_sourceRegister ? registerTagMap_5_valid : _GEN_1526; // @[ReorderBuffer.scala 155:{41,41}]
  wire  _GEN_1528 = 5'h6 == io_decoders_0_source1_sourceRegister ? registerTagMap_6_valid : _GEN_1527; // @[ReorderBuffer.scala 155:{41,41}]
  wire  _GEN_1529 = 5'h7 == io_decoders_0_source1_sourceRegister ? registerTagMap_7_valid : _GEN_1528; // @[ReorderBuffer.scala 155:{41,41}]
  wire  _GEN_1530 = 5'h8 == io_decoders_0_source1_sourceRegister ? registerTagMap_8_valid : _GEN_1529; // @[ReorderBuffer.scala 155:{41,41}]
  wire  _GEN_1531 = 5'h9 == io_decoders_0_source1_sourceRegister ? registerTagMap_9_valid : _GEN_1530; // @[ReorderBuffer.scala 155:{41,41}]
  wire  _GEN_1532 = 5'ha == io_decoders_0_source1_sourceRegister ? registerTagMap_10_valid : _GEN_1531; // @[ReorderBuffer.scala 155:{41,41}]
  wire  _GEN_1533 = 5'hb == io_decoders_0_source1_sourceRegister ? registerTagMap_11_valid : _GEN_1532; // @[ReorderBuffer.scala 155:{41,41}]
  wire  _GEN_1534 = 5'hc == io_decoders_0_source1_sourceRegister ? registerTagMap_12_valid : _GEN_1533; // @[ReorderBuffer.scala 155:{41,41}]
  wire  _GEN_1535 = 5'hd == io_decoders_0_source1_sourceRegister ? registerTagMap_13_valid : _GEN_1534; // @[ReorderBuffer.scala 155:{41,41}]
  wire  _GEN_1536 = 5'he == io_decoders_0_source1_sourceRegister ? registerTagMap_14_valid : _GEN_1535; // @[ReorderBuffer.scala 155:{41,41}]
  wire  _GEN_1537 = 5'hf == io_decoders_0_source1_sourceRegister ? registerTagMap_15_valid : _GEN_1536; // @[ReorderBuffer.scala 155:{41,41}]
  wire  _GEN_1538 = 5'h10 == io_decoders_0_source1_sourceRegister ? registerTagMap_16_valid : _GEN_1537; // @[ReorderBuffer.scala 155:{41,41}]
  wire  _GEN_1539 = 5'h11 == io_decoders_0_source1_sourceRegister ? registerTagMap_17_valid : _GEN_1538; // @[ReorderBuffer.scala 155:{41,41}]
  wire  _GEN_1540 = 5'h12 == io_decoders_0_source1_sourceRegister ? registerTagMap_18_valid : _GEN_1539; // @[ReorderBuffer.scala 155:{41,41}]
  wire  _GEN_1541 = 5'h13 == io_decoders_0_source1_sourceRegister ? registerTagMap_19_valid : _GEN_1540; // @[ReorderBuffer.scala 155:{41,41}]
  wire  _GEN_1542 = 5'h14 == io_decoders_0_source1_sourceRegister ? registerTagMap_20_valid : _GEN_1541; // @[ReorderBuffer.scala 155:{41,41}]
  wire  _GEN_1543 = 5'h15 == io_decoders_0_source1_sourceRegister ? registerTagMap_21_valid : _GEN_1542; // @[ReorderBuffer.scala 155:{41,41}]
  wire  _GEN_1544 = 5'h16 == io_decoders_0_source1_sourceRegister ? registerTagMap_22_valid : _GEN_1543; // @[ReorderBuffer.scala 155:{41,41}]
  wire  _GEN_1545 = 5'h17 == io_decoders_0_source1_sourceRegister ? registerTagMap_23_valid : _GEN_1544; // @[ReorderBuffer.scala 155:{41,41}]
  wire  _GEN_1546 = 5'h18 == io_decoders_0_source1_sourceRegister ? registerTagMap_24_valid : _GEN_1545; // @[ReorderBuffer.scala 155:{41,41}]
  wire  _GEN_1547 = 5'h19 == io_decoders_0_source1_sourceRegister ? registerTagMap_25_valid : _GEN_1546; // @[ReorderBuffer.scala 155:{41,41}]
  wire  _GEN_1548 = 5'h1a == io_decoders_0_source1_sourceRegister ? registerTagMap_26_valid : _GEN_1547; // @[ReorderBuffer.scala 155:{41,41}]
  wire  _GEN_1549 = 5'h1b == io_decoders_0_source1_sourceRegister ? registerTagMap_27_valid : _GEN_1548; // @[ReorderBuffer.scala 155:{41,41}]
  wire  _GEN_1550 = 5'h1c == io_decoders_0_source1_sourceRegister ? registerTagMap_28_valid : _GEN_1549; // @[ReorderBuffer.scala 155:{41,41}]
  wire  _GEN_1551 = 5'h1d == io_decoders_0_source1_sourceRegister ? registerTagMap_29_valid : _GEN_1550; // @[ReorderBuffer.scala 155:{41,41}]
  wire  _GEN_1552 = 5'h1e == io_decoders_0_source1_sourceRegister ? registerTagMap_30_valid : _GEN_1551; // @[ReorderBuffer.scala 155:{41,41}]
  wire  _GEN_1553 = 5'h1f == io_decoders_0_source1_sourceRegister ? registerTagMap_31_valid : _GEN_1552; // @[ReorderBuffer.scala 155:{41,41}]
  wire [3:0] _GEN_1555 = 5'h1 == io_decoders_0_source1_sourceRegister ? registerTagMap_1_tagId : 4'h0; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1556 = 5'h2 == io_decoders_0_source1_sourceRegister ? registerTagMap_2_tagId : _GEN_1555; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1557 = 5'h3 == io_decoders_0_source1_sourceRegister ? registerTagMap_3_tagId : _GEN_1556; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1558 = 5'h4 == io_decoders_0_source1_sourceRegister ? registerTagMap_4_tagId : _GEN_1557; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1559 = 5'h5 == io_decoders_0_source1_sourceRegister ? registerTagMap_5_tagId : _GEN_1558; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1560 = 5'h6 == io_decoders_0_source1_sourceRegister ? registerTagMap_6_tagId : _GEN_1559; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1561 = 5'h7 == io_decoders_0_source1_sourceRegister ? registerTagMap_7_tagId : _GEN_1560; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1562 = 5'h8 == io_decoders_0_source1_sourceRegister ? registerTagMap_8_tagId : _GEN_1561; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1563 = 5'h9 == io_decoders_0_source1_sourceRegister ? registerTagMap_9_tagId : _GEN_1562; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1564 = 5'ha == io_decoders_0_source1_sourceRegister ? registerTagMap_10_tagId : _GEN_1563; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1565 = 5'hb == io_decoders_0_source1_sourceRegister ? registerTagMap_11_tagId : _GEN_1564; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1566 = 5'hc == io_decoders_0_source1_sourceRegister ? registerTagMap_12_tagId : _GEN_1565; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1567 = 5'hd == io_decoders_0_source1_sourceRegister ? registerTagMap_13_tagId : _GEN_1566; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1568 = 5'he == io_decoders_0_source1_sourceRegister ? registerTagMap_14_tagId : _GEN_1567; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1569 = 5'hf == io_decoders_0_source1_sourceRegister ? registerTagMap_15_tagId : _GEN_1568; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1570 = 5'h10 == io_decoders_0_source1_sourceRegister ? registerTagMap_16_tagId : _GEN_1569; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1571 = 5'h11 == io_decoders_0_source1_sourceRegister ? registerTagMap_17_tagId : _GEN_1570; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1572 = 5'h12 == io_decoders_0_source1_sourceRegister ? registerTagMap_18_tagId : _GEN_1571; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1573 = 5'h13 == io_decoders_0_source1_sourceRegister ? registerTagMap_19_tagId : _GEN_1572; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1574 = 5'h14 == io_decoders_0_source1_sourceRegister ? registerTagMap_20_tagId : _GEN_1573; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1575 = 5'h15 == io_decoders_0_source1_sourceRegister ? registerTagMap_21_tagId : _GEN_1574; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1576 = 5'h16 == io_decoders_0_source1_sourceRegister ? registerTagMap_22_tagId : _GEN_1575; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1577 = 5'h17 == io_decoders_0_source1_sourceRegister ? registerTagMap_23_tagId : _GEN_1576; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1578 = 5'h18 == io_decoders_0_source1_sourceRegister ? registerTagMap_24_tagId : _GEN_1577; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1579 = 5'h19 == io_decoders_0_source1_sourceRegister ? registerTagMap_25_tagId : _GEN_1578; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1580 = 5'h1a == io_decoders_0_source1_sourceRegister ? registerTagMap_26_tagId : _GEN_1579; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1581 = 5'h1b == io_decoders_0_source1_sourceRegister ? registerTagMap_27_tagId : _GEN_1580; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1582 = 5'h1c == io_decoders_0_source1_sourceRegister ? registerTagMap_28_tagId : _GEN_1581; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1583 = 5'h1d == io_decoders_0_source1_sourceRegister ? registerTagMap_29_tagId : _GEN_1582; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1584 = 5'h1e == io_decoders_0_source1_sourceRegister ? registerTagMap_30_tagId : _GEN_1583; // @[Tag.scala 23:{10,10}]
  wire [3:0] io_decoders_0_source1_matchingTag_bits_w_id = 5'h1f == io_decoders_0_source1_sourceRegister ?
    registerTagMap_31_tagId : _GEN_1584; // @[Tag.scala 23:{10,10}]
  wire  _GEN_1587 = 4'h1 == io_decoders_0_source1_matchingTag_bits_w_id ? buffer_1_valueReady : buffer_0_valueReady; // @[ReorderBuffer.scala 160:{35,35}]
  wire  _GEN_1588 = 4'h2 == io_decoders_0_source1_matchingTag_bits_w_id ? buffer_2_valueReady : _GEN_1587; // @[ReorderBuffer.scala 160:{35,35}]
  wire  _GEN_1589 = 4'h3 == io_decoders_0_source1_matchingTag_bits_w_id ? buffer_3_valueReady : _GEN_1588; // @[ReorderBuffer.scala 160:{35,35}]
  wire  _GEN_1590 = 4'h4 == io_decoders_0_source1_matchingTag_bits_w_id ? buffer_4_valueReady : _GEN_1589; // @[ReorderBuffer.scala 160:{35,35}]
  wire  _GEN_1591 = 4'h5 == io_decoders_0_source1_matchingTag_bits_w_id ? buffer_5_valueReady : _GEN_1590; // @[ReorderBuffer.scala 160:{35,35}]
  wire  _GEN_1592 = 4'h6 == io_decoders_0_source1_matchingTag_bits_w_id ? buffer_6_valueReady : _GEN_1591; // @[ReorderBuffer.scala 160:{35,35}]
  wire  _GEN_1593 = 4'h7 == io_decoders_0_source1_matchingTag_bits_w_id ? buffer_7_valueReady : _GEN_1592; // @[ReorderBuffer.scala 160:{35,35}]
  wire  _GEN_1594 = 4'h8 == io_decoders_0_source1_matchingTag_bits_w_id ? buffer_8_valueReady : _GEN_1593; // @[ReorderBuffer.scala 160:{35,35}]
  wire  _GEN_1595 = 4'h9 == io_decoders_0_source1_matchingTag_bits_w_id ? buffer_9_valueReady : _GEN_1594; // @[ReorderBuffer.scala 160:{35,35}]
  wire  _GEN_1596 = 4'ha == io_decoders_0_source1_matchingTag_bits_w_id ? buffer_10_valueReady : _GEN_1595; // @[ReorderBuffer.scala 160:{35,35}]
  wire  _GEN_1597 = 4'hb == io_decoders_0_source1_matchingTag_bits_w_id ? buffer_11_valueReady : _GEN_1596; // @[ReorderBuffer.scala 160:{35,35}]
  wire  _GEN_1598 = 4'hc == io_decoders_0_source1_matchingTag_bits_w_id ? buffer_12_valueReady : _GEN_1597; // @[ReorderBuffer.scala 160:{35,35}]
  wire  _GEN_1599 = 4'hd == io_decoders_0_source1_matchingTag_bits_w_id ? buffer_13_valueReady : _GEN_1598; // @[ReorderBuffer.scala 160:{35,35}]
  wire  _GEN_1600 = 4'he == io_decoders_0_source1_matchingTag_bits_w_id ? buffer_14_valueReady : _GEN_1599; // @[ReorderBuffer.scala 160:{35,35}]
  wire  _GEN_1601 = 4'hf == io_decoders_0_source1_matchingTag_bits_w_id ? buffer_15_valueReady : _GEN_1600; // @[ReorderBuffer.scala 160:{35,35}]
  wire [63:0] _GEN_1603 = 4'h1 == io_decoders_0_source1_matchingTag_bits_w_id ? buffer_1_value : buffer_0_value; // @[ReorderBuffer.scala 161:{34,34}]
  wire [63:0] _GEN_1604 = 4'h2 == io_decoders_0_source1_matchingTag_bits_w_id ? buffer_2_value : _GEN_1603; // @[ReorderBuffer.scala 161:{34,34}]
  wire [63:0] _GEN_1605 = 4'h3 == io_decoders_0_source1_matchingTag_bits_w_id ? buffer_3_value : _GEN_1604; // @[ReorderBuffer.scala 161:{34,34}]
  wire [63:0] _GEN_1606 = 4'h4 == io_decoders_0_source1_matchingTag_bits_w_id ? buffer_4_value : _GEN_1605; // @[ReorderBuffer.scala 161:{34,34}]
  wire [63:0] _GEN_1607 = 4'h5 == io_decoders_0_source1_matchingTag_bits_w_id ? buffer_5_value : _GEN_1606; // @[ReorderBuffer.scala 161:{34,34}]
  wire [63:0] _GEN_1608 = 4'h6 == io_decoders_0_source1_matchingTag_bits_w_id ? buffer_6_value : _GEN_1607; // @[ReorderBuffer.scala 161:{34,34}]
  wire [63:0] _GEN_1609 = 4'h7 == io_decoders_0_source1_matchingTag_bits_w_id ? buffer_7_value : _GEN_1608; // @[ReorderBuffer.scala 161:{34,34}]
  wire [63:0] _GEN_1610 = 4'h8 == io_decoders_0_source1_matchingTag_bits_w_id ? buffer_8_value : _GEN_1609; // @[ReorderBuffer.scala 161:{34,34}]
  wire [63:0] _GEN_1611 = 4'h9 == io_decoders_0_source1_matchingTag_bits_w_id ? buffer_9_value : _GEN_1610; // @[ReorderBuffer.scala 161:{34,34}]
  wire [63:0] _GEN_1612 = 4'ha == io_decoders_0_source1_matchingTag_bits_w_id ? buffer_10_value : _GEN_1611; // @[ReorderBuffer.scala 161:{34,34}]
  wire [63:0] _GEN_1613 = 4'hb == io_decoders_0_source1_matchingTag_bits_w_id ? buffer_11_value : _GEN_1612; // @[ReorderBuffer.scala 161:{34,34}]
  wire [63:0] _GEN_1614 = 4'hc == io_decoders_0_source1_matchingTag_bits_w_id ? buffer_12_value : _GEN_1613; // @[ReorderBuffer.scala 161:{34,34}]
  wire [63:0] _GEN_1615 = 4'hd == io_decoders_0_source1_matchingTag_bits_w_id ? buffer_13_value : _GEN_1614; // @[ReorderBuffer.scala 161:{34,34}]
  wire [63:0] _GEN_1616 = 4'he == io_decoders_0_source1_matchingTag_bits_w_id ? buffer_14_value : _GEN_1615; // @[ReorderBuffer.scala 161:{34,34}]
  wire [63:0] _GEN_1617 = 4'hf == io_decoders_0_source1_matchingTag_bits_w_id ? buffer_15_value : _GEN_1616; // @[ReorderBuffer.scala 161:{34,34}]
  wire  _GEN_1625 = 5'h2 == io_decoders_0_source2_sourceRegister ? registerTagMap_2_valid : 5'h1 ==
    io_decoders_0_source2_sourceRegister & registerTagMap_1_valid; // @[ReorderBuffer.scala 172:{41,41}]
  wire  _GEN_1626 = 5'h3 == io_decoders_0_source2_sourceRegister ? registerTagMap_3_valid : _GEN_1625; // @[ReorderBuffer.scala 172:{41,41}]
  wire  _GEN_1627 = 5'h4 == io_decoders_0_source2_sourceRegister ? registerTagMap_4_valid : _GEN_1626; // @[ReorderBuffer.scala 172:{41,41}]
  wire  _GEN_1628 = 5'h5 == io_decoders_0_source2_sourceRegister ? registerTagMap_5_valid : _GEN_1627; // @[ReorderBuffer.scala 172:{41,41}]
  wire  _GEN_1629 = 5'h6 == io_decoders_0_source2_sourceRegister ? registerTagMap_6_valid : _GEN_1628; // @[ReorderBuffer.scala 172:{41,41}]
  wire  _GEN_1630 = 5'h7 == io_decoders_0_source2_sourceRegister ? registerTagMap_7_valid : _GEN_1629; // @[ReorderBuffer.scala 172:{41,41}]
  wire  _GEN_1631 = 5'h8 == io_decoders_0_source2_sourceRegister ? registerTagMap_8_valid : _GEN_1630; // @[ReorderBuffer.scala 172:{41,41}]
  wire  _GEN_1632 = 5'h9 == io_decoders_0_source2_sourceRegister ? registerTagMap_9_valid : _GEN_1631; // @[ReorderBuffer.scala 172:{41,41}]
  wire  _GEN_1633 = 5'ha == io_decoders_0_source2_sourceRegister ? registerTagMap_10_valid : _GEN_1632; // @[ReorderBuffer.scala 172:{41,41}]
  wire  _GEN_1634 = 5'hb == io_decoders_0_source2_sourceRegister ? registerTagMap_11_valid : _GEN_1633; // @[ReorderBuffer.scala 172:{41,41}]
  wire  _GEN_1635 = 5'hc == io_decoders_0_source2_sourceRegister ? registerTagMap_12_valid : _GEN_1634; // @[ReorderBuffer.scala 172:{41,41}]
  wire  _GEN_1636 = 5'hd == io_decoders_0_source2_sourceRegister ? registerTagMap_13_valid : _GEN_1635; // @[ReorderBuffer.scala 172:{41,41}]
  wire  _GEN_1637 = 5'he == io_decoders_0_source2_sourceRegister ? registerTagMap_14_valid : _GEN_1636; // @[ReorderBuffer.scala 172:{41,41}]
  wire  _GEN_1638 = 5'hf == io_decoders_0_source2_sourceRegister ? registerTagMap_15_valid : _GEN_1637; // @[ReorderBuffer.scala 172:{41,41}]
  wire  _GEN_1639 = 5'h10 == io_decoders_0_source2_sourceRegister ? registerTagMap_16_valid : _GEN_1638; // @[ReorderBuffer.scala 172:{41,41}]
  wire  _GEN_1640 = 5'h11 == io_decoders_0_source2_sourceRegister ? registerTagMap_17_valid : _GEN_1639; // @[ReorderBuffer.scala 172:{41,41}]
  wire  _GEN_1641 = 5'h12 == io_decoders_0_source2_sourceRegister ? registerTagMap_18_valid : _GEN_1640; // @[ReorderBuffer.scala 172:{41,41}]
  wire  _GEN_1642 = 5'h13 == io_decoders_0_source2_sourceRegister ? registerTagMap_19_valid : _GEN_1641; // @[ReorderBuffer.scala 172:{41,41}]
  wire  _GEN_1643 = 5'h14 == io_decoders_0_source2_sourceRegister ? registerTagMap_20_valid : _GEN_1642; // @[ReorderBuffer.scala 172:{41,41}]
  wire  _GEN_1644 = 5'h15 == io_decoders_0_source2_sourceRegister ? registerTagMap_21_valid : _GEN_1643; // @[ReorderBuffer.scala 172:{41,41}]
  wire  _GEN_1645 = 5'h16 == io_decoders_0_source2_sourceRegister ? registerTagMap_22_valid : _GEN_1644; // @[ReorderBuffer.scala 172:{41,41}]
  wire  _GEN_1646 = 5'h17 == io_decoders_0_source2_sourceRegister ? registerTagMap_23_valid : _GEN_1645; // @[ReorderBuffer.scala 172:{41,41}]
  wire  _GEN_1647 = 5'h18 == io_decoders_0_source2_sourceRegister ? registerTagMap_24_valid : _GEN_1646; // @[ReorderBuffer.scala 172:{41,41}]
  wire  _GEN_1648 = 5'h19 == io_decoders_0_source2_sourceRegister ? registerTagMap_25_valid : _GEN_1647; // @[ReorderBuffer.scala 172:{41,41}]
  wire  _GEN_1649 = 5'h1a == io_decoders_0_source2_sourceRegister ? registerTagMap_26_valid : _GEN_1648; // @[ReorderBuffer.scala 172:{41,41}]
  wire  _GEN_1650 = 5'h1b == io_decoders_0_source2_sourceRegister ? registerTagMap_27_valid : _GEN_1649; // @[ReorderBuffer.scala 172:{41,41}]
  wire  _GEN_1651 = 5'h1c == io_decoders_0_source2_sourceRegister ? registerTagMap_28_valid : _GEN_1650; // @[ReorderBuffer.scala 172:{41,41}]
  wire  _GEN_1652 = 5'h1d == io_decoders_0_source2_sourceRegister ? registerTagMap_29_valid : _GEN_1651; // @[ReorderBuffer.scala 172:{41,41}]
  wire  _GEN_1653 = 5'h1e == io_decoders_0_source2_sourceRegister ? registerTagMap_30_valid : _GEN_1652; // @[ReorderBuffer.scala 172:{41,41}]
  wire  _GEN_1654 = 5'h1f == io_decoders_0_source2_sourceRegister ? registerTagMap_31_valid : _GEN_1653; // @[ReorderBuffer.scala 172:{41,41}]
  wire [3:0] _GEN_1656 = 5'h1 == io_decoders_0_source2_sourceRegister ? registerTagMap_1_tagId : 4'h0; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1657 = 5'h2 == io_decoders_0_source2_sourceRegister ? registerTagMap_2_tagId : _GEN_1656; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1658 = 5'h3 == io_decoders_0_source2_sourceRegister ? registerTagMap_3_tagId : _GEN_1657; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1659 = 5'h4 == io_decoders_0_source2_sourceRegister ? registerTagMap_4_tagId : _GEN_1658; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1660 = 5'h5 == io_decoders_0_source2_sourceRegister ? registerTagMap_5_tagId : _GEN_1659; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1661 = 5'h6 == io_decoders_0_source2_sourceRegister ? registerTagMap_6_tagId : _GEN_1660; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1662 = 5'h7 == io_decoders_0_source2_sourceRegister ? registerTagMap_7_tagId : _GEN_1661; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1663 = 5'h8 == io_decoders_0_source2_sourceRegister ? registerTagMap_8_tagId : _GEN_1662; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1664 = 5'h9 == io_decoders_0_source2_sourceRegister ? registerTagMap_9_tagId : _GEN_1663; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1665 = 5'ha == io_decoders_0_source2_sourceRegister ? registerTagMap_10_tagId : _GEN_1664; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1666 = 5'hb == io_decoders_0_source2_sourceRegister ? registerTagMap_11_tagId : _GEN_1665; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1667 = 5'hc == io_decoders_0_source2_sourceRegister ? registerTagMap_12_tagId : _GEN_1666; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1668 = 5'hd == io_decoders_0_source2_sourceRegister ? registerTagMap_13_tagId : _GEN_1667; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1669 = 5'he == io_decoders_0_source2_sourceRegister ? registerTagMap_14_tagId : _GEN_1668; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1670 = 5'hf == io_decoders_0_source2_sourceRegister ? registerTagMap_15_tagId : _GEN_1669; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1671 = 5'h10 == io_decoders_0_source2_sourceRegister ? registerTagMap_16_tagId : _GEN_1670; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1672 = 5'h11 == io_decoders_0_source2_sourceRegister ? registerTagMap_17_tagId : _GEN_1671; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1673 = 5'h12 == io_decoders_0_source2_sourceRegister ? registerTagMap_18_tagId : _GEN_1672; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1674 = 5'h13 == io_decoders_0_source2_sourceRegister ? registerTagMap_19_tagId : _GEN_1673; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1675 = 5'h14 == io_decoders_0_source2_sourceRegister ? registerTagMap_20_tagId : _GEN_1674; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1676 = 5'h15 == io_decoders_0_source2_sourceRegister ? registerTagMap_21_tagId : _GEN_1675; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1677 = 5'h16 == io_decoders_0_source2_sourceRegister ? registerTagMap_22_tagId : _GEN_1676; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1678 = 5'h17 == io_decoders_0_source2_sourceRegister ? registerTagMap_23_tagId : _GEN_1677; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1679 = 5'h18 == io_decoders_0_source2_sourceRegister ? registerTagMap_24_tagId : _GEN_1678; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1680 = 5'h19 == io_decoders_0_source2_sourceRegister ? registerTagMap_25_tagId : _GEN_1679; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1681 = 5'h1a == io_decoders_0_source2_sourceRegister ? registerTagMap_26_tagId : _GEN_1680; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1682 = 5'h1b == io_decoders_0_source2_sourceRegister ? registerTagMap_27_tagId : _GEN_1681; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1683 = 5'h1c == io_decoders_0_source2_sourceRegister ? registerTagMap_28_tagId : _GEN_1682; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1684 = 5'h1d == io_decoders_0_source2_sourceRegister ? registerTagMap_29_tagId : _GEN_1683; // @[Tag.scala 23:{10,10}]
  wire [3:0] _GEN_1685 = 5'h1e == io_decoders_0_source2_sourceRegister ? registerTagMap_30_tagId : _GEN_1684; // @[Tag.scala 23:{10,10}]
  wire [3:0] io_decoders_0_source2_matchingTag_bits_w_id = 5'h1f == io_decoders_0_source2_sourceRegister ?
    registerTagMap_31_tagId : _GEN_1685; // @[Tag.scala 23:{10,10}]
  wire  _GEN_1688 = 4'h1 == io_decoders_0_source2_matchingTag_bits_w_id ? buffer_1_valueReady : buffer_0_valueReady; // @[ReorderBuffer.scala 177:{35,35}]
  wire  _GEN_1689 = 4'h2 == io_decoders_0_source2_matchingTag_bits_w_id ? buffer_2_valueReady : _GEN_1688; // @[ReorderBuffer.scala 177:{35,35}]
  wire  _GEN_1690 = 4'h3 == io_decoders_0_source2_matchingTag_bits_w_id ? buffer_3_valueReady : _GEN_1689; // @[ReorderBuffer.scala 177:{35,35}]
  wire  _GEN_1691 = 4'h4 == io_decoders_0_source2_matchingTag_bits_w_id ? buffer_4_valueReady : _GEN_1690; // @[ReorderBuffer.scala 177:{35,35}]
  wire  _GEN_1692 = 4'h5 == io_decoders_0_source2_matchingTag_bits_w_id ? buffer_5_valueReady : _GEN_1691; // @[ReorderBuffer.scala 177:{35,35}]
  wire  _GEN_1693 = 4'h6 == io_decoders_0_source2_matchingTag_bits_w_id ? buffer_6_valueReady : _GEN_1692; // @[ReorderBuffer.scala 177:{35,35}]
  wire  _GEN_1694 = 4'h7 == io_decoders_0_source2_matchingTag_bits_w_id ? buffer_7_valueReady : _GEN_1693; // @[ReorderBuffer.scala 177:{35,35}]
  wire  _GEN_1695 = 4'h8 == io_decoders_0_source2_matchingTag_bits_w_id ? buffer_8_valueReady : _GEN_1694; // @[ReorderBuffer.scala 177:{35,35}]
  wire  _GEN_1696 = 4'h9 == io_decoders_0_source2_matchingTag_bits_w_id ? buffer_9_valueReady : _GEN_1695; // @[ReorderBuffer.scala 177:{35,35}]
  wire  _GEN_1697 = 4'ha == io_decoders_0_source2_matchingTag_bits_w_id ? buffer_10_valueReady : _GEN_1696; // @[ReorderBuffer.scala 177:{35,35}]
  wire  _GEN_1698 = 4'hb == io_decoders_0_source2_matchingTag_bits_w_id ? buffer_11_valueReady : _GEN_1697; // @[ReorderBuffer.scala 177:{35,35}]
  wire  _GEN_1699 = 4'hc == io_decoders_0_source2_matchingTag_bits_w_id ? buffer_12_valueReady : _GEN_1698; // @[ReorderBuffer.scala 177:{35,35}]
  wire  _GEN_1700 = 4'hd == io_decoders_0_source2_matchingTag_bits_w_id ? buffer_13_valueReady : _GEN_1699; // @[ReorderBuffer.scala 177:{35,35}]
  wire  _GEN_1701 = 4'he == io_decoders_0_source2_matchingTag_bits_w_id ? buffer_14_valueReady : _GEN_1700; // @[ReorderBuffer.scala 177:{35,35}]
  wire  _GEN_1702 = 4'hf == io_decoders_0_source2_matchingTag_bits_w_id ? buffer_15_valueReady : _GEN_1701; // @[ReorderBuffer.scala 177:{35,35}]
  wire [63:0] _GEN_1704 = 4'h1 == io_decoders_0_source2_matchingTag_bits_w_id ? buffer_1_value : buffer_0_value; // @[ReorderBuffer.scala 178:{34,34}]
  wire [63:0] _GEN_1705 = 4'h2 == io_decoders_0_source2_matchingTag_bits_w_id ? buffer_2_value : _GEN_1704; // @[ReorderBuffer.scala 178:{34,34}]
  wire [63:0] _GEN_1706 = 4'h3 == io_decoders_0_source2_matchingTag_bits_w_id ? buffer_3_value : _GEN_1705; // @[ReorderBuffer.scala 178:{34,34}]
  wire [63:0] _GEN_1707 = 4'h4 == io_decoders_0_source2_matchingTag_bits_w_id ? buffer_4_value : _GEN_1706; // @[ReorderBuffer.scala 178:{34,34}]
  wire [63:0] _GEN_1708 = 4'h5 == io_decoders_0_source2_matchingTag_bits_w_id ? buffer_5_value : _GEN_1707; // @[ReorderBuffer.scala 178:{34,34}]
  wire [63:0] _GEN_1709 = 4'h6 == io_decoders_0_source2_matchingTag_bits_w_id ? buffer_6_value : _GEN_1708; // @[ReorderBuffer.scala 178:{34,34}]
  wire [63:0] _GEN_1710 = 4'h7 == io_decoders_0_source2_matchingTag_bits_w_id ? buffer_7_value : _GEN_1709; // @[ReorderBuffer.scala 178:{34,34}]
  wire [63:0] _GEN_1711 = 4'h8 == io_decoders_0_source2_matchingTag_bits_w_id ? buffer_8_value : _GEN_1710; // @[ReorderBuffer.scala 178:{34,34}]
  wire [63:0] _GEN_1712 = 4'h9 == io_decoders_0_source2_matchingTag_bits_w_id ? buffer_9_value : _GEN_1711; // @[ReorderBuffer.scala 178:{34,34}]
  wire [63:0] _GEN_1713 = 4'ha == io_decoders_0_source2_matchingTag_bits_w_id ? buffer_10_value : _GEN_1712; // @[ReorderBuffer.scala 178:{34,34}]
  wire [63:0] _GEN_1714 = 4'hb == io_decoders_0_source2_matchingTag_bits_w_id ? buffer_11_value : _GEN_1713; // @[ReorderBuffer.scala 178:{34,34}]
  wire [63:0] _GEN_1715 = 4'hc == io_decoders_0_source2_matchingTag_bits_w_id ? buffer_12_value : _GEN_1714; // @[ReorderBuffer.scala 178:{34,34}]
  wire [63:0] _GEN_1716 = 4'hd == io_decoders_0_source2_matchingTag_bits_w_id ? buffer_13_value : _GEN_1715; // @[ReorderBuffer.scala 178:{34,34}]
  wire [63:0] _GEN_1717 = 4'he == io_decoders_0_source2_matchingTag_bits_w_id ? buffer_14_value : _GEN_1716; // @[ReorderBuffer.scala 178:{34,34}]
  wire [63:0] _GEN_1718 = 4'hf == io_decoders_0_source2_matchingTag_bits_w_id ? buffer_15_value : _GEN_1717; // @[ReorderBuffer.scala 178:{34,34}]
  wire [3:0] _GEN_1853 = {{1'd0}, tailDelta}; // @[ReorderBuffer.scala 193:45]
  wire [3:0] _tail_T_1 = tail + _GEN_1853; // @[ReorderBuffer.scala 193:45]
  wire [2:0] _io_csr_retireCount_T = io_isError ? 3'h0 : tailDelta; // @[ReorderBuffer.scala 194:28]
  wire  _T_19 = io_collectedOutputs_outputs_valid & ~io_collectedOutputs_outputs_bits_resultType &
    io_collectedOutputs_outputs_bits_tag_threadId; // @[ReorderBuffer.scala 200:68]
  wire  _GEN_1756 = 4'h0 == io_collectedOutputs_outputs_bits_tag_id | _GEN_1314; // @[ReorderBuffer.scala 204:{43,43}]
  wire  _GEN_1757 = 4'h1 == io_collectedOutputs_outputs_bits_tag_id | _GEN_1315; // @[ReorderBuffer.scala 204:{43,43}]
  wire  _GEN_1758 = 4'h2 == io_collectedOutputs_outputs_bits_tag_id | _GEN_1316; // @[ReorderBuffer.scala 204:{43,43}]
  wire  _GEN_1759 = 4'h3 == io_collectedOutputs_outputs_bits_tag_id | _GEN_1317; // @[ReorderBuffer.scala 204:{43,43}]
  wire  _GEN_1760 = 4'h4 == io_collectedOutputs_outputs_bits_tag_id | _GEN_1318; // @[ReorderBuffer.scala 204:{43,43}]
  wire  _GEN_1761 = 4'h5 == io_collectedOutputs_outputs_bits_tag_id | _GEN_1319; // @[ReorderBuffer.scala 204:{43,43}]
  wire  _GEN_1762 = 4'h6 == io_collectedOutputs_outputs_bits_tag_id | _GEN_1320; // @[ReorderBuffer.scala 204:{43,43}]
  wire  _GEN_1763 = 4'h7 == io_collectedOutputs_outputs_bits_tag_id | _GEN_1321; // @[ReorderBuffer.scala 204:{43,43}]
  wire  _GEN_1764 = 4'h8 == io_collectedOutputs_outputs_bits_tag_id | _GEN_1322; // @[ReorderBuffer.scala 204:{43,43}]
  wire  _GEN_1765 = 4'h9 == io_collectedOutputs_outputs_bits_tag_id | _GEN_1323; // @[ReorderBuffer.scala 204:{43,43}]
  wire  _GEN_1766 = 4'ha == io_collectedOutputs_outputs_bits_tag_id | _GEN_1324; // @[ReorderBuffer.scala 204:{43,43}]
  wire  _GEN_1767 = 4'hb == io_collectedOutputs_outputs_bits_tag_id | _GEN_1325; // @[ReorderBuffer.scala 204:{43,43}]
  wire  _GEN_1768 = 4'hc == io_collectedOutputs_outputs_bits_tag_id | _GEN_1326; // @[ReorderBuffer.scala 204:{43,43}]
  wire  _GEN_1769 = 4'hd == io_collectedOutputs_outputs_bits_tag_id | _GEN_1327; // @[ReorderBuffer.scala 204:{43,43}]
  wire  _GEN_1770 = 4'he == io_collectedOutputs_outputs_bits_tag_id | _GEN_1328; // @[ReorderBuffer.scala 204:{43,43}]
  wire  _GEN_1771 = 4'hf == io_collectedOutputs_outputs_bits_tag_id | _GEN_1329; // @[ReorderBuffer.scala 204:{43,43}]
  assign io_decoders_0_source1_matchingTag_valid = io_decoders_0_source1_sourceRegister != 5'h0 & _GEN_1553; // @[ReorderBuffer.scala 151:50 155:41 163:41]
  assign io_decoders_0_source1_matchingTag_bits_id = io_decoders_0_source1_sourceRegister != 5'h0 ?
    io_decoders_0_source1_matchingTag_bits_w_id : 4'h0; // @[ReorderBuffer.scala 151:50 156:40 164:40]
  assign io_decoders_0_source1_value_valid = io_decoders_0_source1_sourceRegister != 5'h0 & _GEN_1601; // @[ReorderBuffer.scala 151:50 160:35 165:35]
  assign io_decoders_0_source1_value_bits = io_decoders_0_source1_sourceRegister != 5'h0 ? _GEN_1617 : 64'h0; // @[ReorderBuffer.scala 151:50 161:34 166:34]
  assign io_decoders_0_source2_matchingTag_valid = io_decoders_0_source2_sourceRegister != 5'h0 & _GEN_1654; // @[ReorderBuffer.scala 169:50 172:41 180:41]
  assign io_decoders_0_source2_matchingTag_bits_id = io_decoders_0_source2_sourceRegister != 5'h0 ?
    io_decoders_0_source2_matchingTag_bits_w_id : 4'h0; // @[ReorderBuffer.scala 169:50 173:40 181:40]
  assign io_decoders_0_source2_value_valid = io_decoders_0_source2_sourceRegister != 5'h0 & _GEN_1702; // @[ReorderBuffer.scala 169:50 177:35 182:35]
  assign io_decoders_0_source2_value_bits = io_decoders_0_source2_sourceRegister != 5'h0 ? _GEN_1718 : 64'h0; // @[ReorderBuffer.scala 169:50 178:34 183:34]
  assign io_decoders_0_destination_destinationTag_id = head; // @[Tag.scala 21:17 23:10]
  assign io_decoders_0_ready = _io_decoders_0_ready_T_1 != tail; // @[ReorderBuffer.scala 129:55]
  assign io_registerFile_0_valid = canCommit & ~_GEN_47; // @[ReorderBuffer.scala 83:27]
  assign io_registerFile_0_bits_destinationRegister = canCommit ? _GEN_209 : 5'h0; // @[ReorderBuffer.scala 88:21 85:33]
  assign io_registerFile_0_bits_value = canCommit ? _GEN_208 : 64'h0; // @[ReorderBuffer.scala 84:19 88:21]
  assign io_registerFile_1_valid = canCommit_1 & ~_GEN_346; // @[ReorderBuffer.scala 83:27]
  assign io_registerFile_1_bits_destinationRegister = canCommit_1 ? _GEN_508 : 5'h0; // @[ReorderBuffer.scala 88:21 85:33]
  assign io_registerFile_1_bits_value = canCommit_1 ? _GEN_507 : 64'h0; // @[ReorderBuffer.scala 84:19 88:21]
  assign io_registerFile_2_valid = canCommit_2 & ~_GEN_647; // @[ReorderBuffer.scala 83:27]
  assign io_registerFile_2_bits_destinationRegister = canCommit_2 ? _GEN_809 : 5'h0; // @[ReorderBuffer.scala 88:21 85:33]
  assign io_registerFile_2_bits_value = canCommit_2 ? _GEN_808 : 64'h0; // @[ReorderBuffer.scala 84:19 88:21]
  assign io_registerFile_3_valid = canCommit_3 & ~_GEN_948; // @[ReorderBuffer.scala 83:27]
  assign io_registerFile_3_bits_destinationRegister = canCommit_3 ? _GEN_1110 : 5'h0; // @[ReorderBuffer.scala 88:21 85:33]
  assign io_registerFile_3_bits_value = canCommit_3 ? _GEN_1109 : 64'h0; // @[ReorderBuffer.scala 84:19 88:21]
  assign io_loadStoreQueue_0_valid = canCommit & _GEN_31; // @[ReorderBuffer.scala 106:21 109:17 113:17]
  assign io_loadStoreQueue_0_bits_destinationTag_id = canCommit ? index : 4'h0; // @[ReorderBuffer.scala 106:21 108:31 112:31]
  assign io_loadStoreQueue_1_valid = canCommit_1 & _GEN_330; // @[ReorderBuffer.scala 106:21 109:17 113:17]
  assign io_loadStoreQueue_1_bits_destinationTag_id = canCommit_1 ? index_1 : 4'h0; // @[ReorderBuffer.scala 106:21 108:31 112:31]
  assign io_loadStoreQueue_2_valid = canCommit_2 & _GEN_631; // @[ReorderBuffer.scala 106:21 109:17 113:17]
  assign io_loadStoreQueue_2_bits_destinationTag_id = canCommit_2 ? index_2 : 4'h0; // @[ReorderBuffer.scala 106:21 108:31 112:31]
  assign io_loadStoreQueue_3_valid = canCommit_3 & _GEN_932; // @[ReorderBuffer.scala 106:21 109:17 113:17]
  assign io_loadStoreQueue_3_bits_destinationTag_id = canCommit_3 ? index_3 : 4'h0; // @[ReorderBuffer.scala 106:21 108:31 112:31]
  assign io_isEmpty = head == tail; // @[ReorderBuffer.scala 195:22]
  assign io_csr_retireCount = _io_csr_retireCount_T[1:0]; // @[ReorderBuffer.scala 194:22]
  assign io_isError = canCommit_3 ? _GEN_1145 : _GEN_881; // @[ReorderBuffer.scala 88:21]
  always @(posedge clock) begin
    if (reset) begin // @[ReorderBuffer.scala 53:21]
      head <= 4'h0; // @[ReorderBuffer.scala 53:21]
    end else if (_T_8) begin // @[ReorderBuffer.scala 189:10]
      head <= _io_decoders_0_ready_T_1;
    end
    if (reset) begin // @[ReorderBuffer.scala 54:21]
      tail <= 4'h0; // @[ReorderBuffer.scala 54:21]
    end else if (io_isError) begin // @[ReorderBuffer.scala 193:14]
      if (_T_8) begin // @[ReorderBuffer.scala 189:10]
        tail <= _io_decoders_0_ready_T_1;
      end else begin
        tail <= head;
      end
    end else begin
      tail <= _tail_T_1;
    end
    if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'h0 == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_0_destinationRegister <= io_decoders_0_destination_destinationRegister; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      buffer_0_valueReady <= _GEN_1756;
    end else if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'h0 == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_0_valueReady <= 1'h0; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      if (4'h0 == io_collectedOutputs_outputs_bits_tag_id) begin // @[ReorderBuffer.scala 202:38]
        buffer_0_value <= io_collectedOutputs_outputs_bits_value; // @[ReorderBuffer.scala 202:38]
      end else begin
        buffer_0_value <= _GEN_1330;
      end
    end else begin
      buffer_0_value <= _GEN_1330;
    end
    if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'h0 == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_0_storeSign <= io_decoders_0_destination_storeSign; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      if (4'h0 == io_collectedOutputs_outputs_bits_tag_id) begin // @[ReorderBuffer.scala 203:40]
        buffer_0_isError <= io_collectedOutputs_outputs_bits_isError; // @[ReorderBuffer.scala 203:40]
      end else begin
        buffer_0_isError <= _GEN_1378;
      end
    end else begin
      buffer_0_isError <= _GEN_1378;
    end
    if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'h1 == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_1_destinationRegister <= io_decoders_0_destination_destinationRegister; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      buffer_1_valueReady <= _GEN_1757;
    end else if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'h1 == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_1_valueReady <= 1'h0; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      if (4'h1 == io_collectedOutputs_outputs_bits_tag_id) begin // @[ReorderBuffer.scala 202:38]
        buffer_1_value <= io_collectedOutputs_outputs_bits_value; // @[ReorderBuffer.scala 202:38]
      end else begin
        buffer_1_value <= _GEN_1331;
      end
    end else begin
      buffer_1_value <= _GEN_1331;
    end
    if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'h1 == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_1_storeSign <= io_decoders_0_destination_storeSign; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      if (4'h1 == io_collectedOutputs_outputs_bits_tag_id) begin // @[ReorderBuffer.scala 203:40]
        buffer_1_isError <= io_collectedOutputs_outputs_bits_isError; // @[ReorderBuffer.scala 203:40]
      end else begin
        buffer_1_isError <= _GEN_1379;
      end
    end else begin
      buffer_1_isError <= _GEN_1379;
    end
    if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'h2 == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_2_destinationRegister <= io_decoders_0_destination_destinationRegister; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      buffer_2_valueReady <= _GEN_1758;
    end else if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'h2 == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_2_valueReady <= 1'h0; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      if (4'h2 == io_collectedOutputs_outputs_bits_tag_id) begin // @[ReorderBuffer.scala 202:38]
        buffer_2_value <= io_collectedOutputs_outputs_bits_value; // @[ReorderBuffer.scala 202:38]
      end else begin
        buffer_2_value <= _GEN_1332;
      end
    end else begin
      buffer_2_value <= _GEN_1332;
    end
    if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'h2 == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_2_storeSign <= io_decoders_0_destination_storeSign; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      if (4'h2 == io_collectedOutputs_outputs_bits_tag_id) begin // @[ReorderBuffer.scala 203:40]
        buffer_2_isError <= io_collectedOutputs_outputs_bits_isError; // @[ReorderBuffer.scala 203:40]
      end else begin
        buffer_2_isError <= _GEN_1380;
      end
    end else begin
      buffer_2_isError <= _GEN_1380;
    end
    if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'h3 == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_3_destinationRegister <= io_decoders_0_destination_destinationRegister; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      buffer_3_valueReady <= _GEN_1759;
    end else if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'h3 == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_3_valueReady <= 1'h0; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      if (4'h3 == io_collectedOutputs_outputs_bits_tag_id) begin // @[ReorderBuffer.scala 202:38]
        buffer_3_value <= io_collectedOutputs_outputs_bits_value; // @[ReorderBuffer.scala 202:38]
      end else begin
        buffer_3_value <= _GEN_1333;
      end
    end else begin
      buffer_3_value <= _GEN_1333;
    end
    if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'h3 == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_3_storeSign <= io_decoders_0_destination_storeSign; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      if (4'h3 == io_collectedOutputs_outputs_bits_tag_id) begin // @[ReorderBuffer.scala 203:40]
        buffer_3_isError <= io_collectedOutputs_outputs_bits_isError; // @[ReorderBuffer.scala 203:40]
      end else begin
        buffer_3_isError <= _GEN_1381;
      end
    end else begin
      buffer_3_isError <= _GEN_1381;
    end
    if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'h4 == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_4_destinationRegister <= io_decoders_0_destination_destinationRegister; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      buffer_4_valueReady <= _GEN_1760;
    end else if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'h4 == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_4_valueReady <= 1'h0; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      if (4'h4 == io_collectedOutputs_outputs_bits_tag_id) begin // @[ReorderBuffer.scala 202:38]
        buffer_4_value <= io_collectedOutputs_outputs_bits_value; // @[ReorderBuffer.scala 202:38]
      end else begin
        buffer_4_value <= _GEN_1334;
      end
    end else begin
      buffer_4_value <= _GEN_1334;
    end
    if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'h4 == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_4_storeSign <= io_decoders_0_destination_storeSign; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      if (4'h4 == io_collectedOutputs_outputs_bits_tag_id) begin // @[ReorderBuffer.scala 203:40]
        buffer_4_isError <= io_collectedOutputs_outputs_bits_isError; // @[ReorderBuffer.scala 203:40]
      end else begin
        buffer_4_isError <= _GEN_1382;
      end
    end else begin
      buffer_4_isError <= _GEN_1382;
    end
    if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'h5 == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_5_destinationRegister <= io_decoders_0_destination_destinationRegister; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      buffer_5_valueReady <= _GEN_1761;
    end else if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'h5 == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_5_valueReady <= 1'h0; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      if (4'h5 == io_collectedOutputs_outputs_bits_tag_id) begin // @[ReorderBuffer.scala 202:38]
        buffer_5_value <= io_collectedOutputs_outputs_bits_value; // @[ReorderBuffer.scala 202:38]
      end else begin
        buffer_5_value <= _GEN_1335;
      end
    end else begin
      buffer_5_value <= _GEN_1335;
    end
    if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'h5 == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_5_storeSign <= io_decoders_0_destination_storeSign; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      if (4'h5 == io_collectedOutputs_outputs_bits_tag_id) begin // @[ReorderBuffer.scala 203:40]
        buffer_5_isError <= io_collectedOutputs_outputs_bits_isError; // @[ReorderBuffer.scala 203:40]
      end else begin
        buffer_5_isError <= _GEN_1383;
      end
    end else begin
      buffer_5_isError <= _GEN_1383;
    end
    if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'h6 == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_6_destinationRegister <= io_decoders_0_destination_destinationRegister; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      buffer_6_valueReady <= _GEN_1762;
    end else if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'h6 == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_6_valueReady <= 1'h0; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      if (4'h6 == io_collectedOutputs_outputs_bits_tag_id) begin // @[ReorderBuffer.scala 202:38]
        buffer_6_value <= io_collectedOutputs_outputs_bits_value; // @[ReorderBuffer.scala 202:38]
      end else begin
        buffer_6_value <= _GEN_1336;
      end
    end else begin
      buffer_6_value <= _GEN_1336;
    end
    if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'h6 == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_6_storeSign <= io_decoders_0_destination_storeSign; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      if (4'h6 == io_collectedOutputs_outputs_bits_tag_id) begin // @[ReorderBuffer.scala 203:40]
        buffer_6_isError <= io_collectedOutputs_outputs_bits_isError; // @[ReorderBuffer.scala 203:40]
      end else begin
        buffer_6_isError <= _GEN_1384;
      end
    end else begin
      buffer_6_isError <= _GEN_1384;
    end
    if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'h7 == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_7_destinationRegister <= io_decoders_0_destination_destinationRegister; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      buffer_7_valueReady <= _GEN_1763;
    end else if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'h7 == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_7_valueReady <= 1'h0; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      if (4'h7 == io_collectedOutputs_outputs_bits_tag_id) begin // @[ReorderBuffer.scala 202:38]
        buffer_7_value <= io_collectedOutputs_outputs_bits_value; // @[ReorderBuffer.scala 202:38]
      end else begin
        buffer_7_value <= _GEN_1337;
      end
    end else begin
      buffer_7_value <= _GEN_1337;
    end
    if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'h7 == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_7_storeSign <= io_decoders_0_destination_storeSign; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      if (4'h7 == io_collectedOutputs_outputs_bits_tag_id) begin // @[ReorderBuffer.scala 203:40]
        buffer_7_isError <= io_collectedOutputs_outputs_bits_isError; // @[ReorderBuffer.scala 203:40]
      end else begin
        buffer_7_isError <= _GEN_1385;
      end
    end else begin
      buffer_7_isError <= _GEN_1385;
    end
    if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'h8 == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_8_destinationRegister <= io_decoders_0_destination_destinationRegister; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      buffer_8_valueReady <= _GEN_1764;
    end else if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'h8 == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_8_valueReady <= 1'h0; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      if (4'h8 == io_collectedOutputs_outputs_bits_tag_id) begin // @[ReorderBuffer.scala 202:38]
        buffer_8_value <= io_collectedOutputs_outputs_bits_value; // @[ReorderBuffer.scala 202:38]
      end else begin
        buffer_8_value <= _GEN_1338;
      end
    end else begin
      buffer_8_value <= _GEN_1338;
    end
    if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'h8 == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_8_storeSign <= io_decoders_0_destination_storeSign; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      if (4'h8 == io_collectedOutputs_outputs_bits_tag_id) begin // @[ReorderBuffer.scala 203:40]
        buffer_8_isError <= io_collectedOutputs_outputs_bits_isError; // @[ReorderBuffer.scala 203:40]
      end else begin
        buffer_8_isError <= _GEN_1386;
      end
    end else begin
      buffer_8_isError <= _GEN_1386;
    end
    if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'h9 == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_9_destinationRegister <= io_decoders_0_destination_destinationRegister; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      buffer_9_valueReady <= _GEN_1765;
    end else if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'h9 == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_9_valueReady <= 1'h0; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      if (4'h9 == io_collectedOutputs_outputs_bits_tag_id) begin // @[ReorderBuffer.scala 202:38]
        buffer_9_value <= io_collectedOutputs_outputs_bits_value; // @[ReorderBuffer.scala 202:38]
      end else begin
        buffer_9_value <= _GEN_1339;
      end
    end else begin
      buffer_9_value <= _GEN_1339;
    end
    if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'h9 == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_9_storeSign <= io_decoders_0_destination_storeSign; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      if (4'h9 == io_collectedOutputs_outputs_bits_tag_id) begin // @[ReorderBuffer.scala 203:40]
        buffer_9_isError <= io_collectedOutputs_outputs_bits_isError; // @[ReorderBuffer.scala 203:40]
      end else begin
        buffer_9_isError <= _GEN_1387;
      end
    end else begin
      buffer_9_isError <= _GEN_1387;
    end
    if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'ha == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_10_destinationRegister <= io_decoders_0_destination_destinationRegister; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      buffer_10_valueReady <= _GEN_1766;
    end else if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'ha == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_10_valueReady <= 1'h0; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      if (4'ha == io_collectedOutputs_outputs_bits_tag_id) begin // @[ReorderBuffer.scala 202:38]
        buffer_10_value <= io_collectedOutputs_outputs_bits_value; // @[ReorderBuffer.scala 202:38]
      end else begin
        buffer_10_value <= _GEN_1340;
      end
    end else begin
      buffer_10_value <= _GEN_1340;
    end
    if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'ha == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_10_storeSign <= io_decoders_0_destination_storeSign; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      if (4'ha == io_collectedOutputs_outputs_bits_tag_id) begin // @[ReorderBuffer.scala 203:40]
        buffer_10_isError <= io_collectedOutputs_outputs_bits_isError; // @[ReorderBuffer.scala 203:40]
      end else begin
        buffer_10_isError <= _GEN_1388;
      end
    end else begin
      buffer_10_isError <= _GEN_1388;
    end
    if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'hb == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_11_destinationRegister <= io_decoders_0_destination_destinationRegister; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      buffer_11_valueReady <= _GEN_1767;
    end else if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'hb == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_11_valueReady <= 1'h0; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      if (4'hb == io_collectedOutputs_outputs_bits_tag_id) begin // @[ReorderBuffer.scala 202:38]
        buffer_11_value <= io_collectedOutputs_outputs_bits_value; // @[ReorderBuffer.scala 202:38]
      end else begin
        buffer_11_value <= _GEN_1341;
      end
    end else begin
      buffer_11_value <= _GEN_1341;
    end
    if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'hb == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_11_storeSign <= io_decoders_0_destination_storeSign; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      if (4'hb == io_collectedOutputs_outputs_bits_tag_id) begin // @[ReorderBuffer.scala 203:40]
        buffer_11_isError <= io_collectedOutputs_outputs_bits_isError; // @[ReorderBuffer.scala 203:40]
      end else begin
        buffer_11_isError <= _GEN_1389;
      end
    end else begin
      buffer_11_isError <= _GEN_1389;
    end
    if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'hc == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_12_destinationRegister <= io_decoders_0_destination_destinationRegister; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      buffer_12_valueReady <= _GEN_1768;
    end else if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'hc == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_12_valueReady <= 1'h0; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      if (4'hc == io_collectedOutputs_outputs_bits_tag_id) begin // @[ReorderBuffer.scala 202:38]
        buffer_12_value <= io_collectedOutputs_outputs_bits_value; // @[ReorderBuffer.scala 202:38]
      end else begin
        buffer_12_value <= _GEN_1342;
      end
    end else begin
      buffer_12_value <= _GEN_1342;
    end
    if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'hc == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_12_storeSign <= io_decoders_0_destination_storeSign; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      if (4'hc == io_collectedOutputs_outputs_bits_tag_id) begin // @[ReorderBuffer.scala 203:40]
        buffer_12_isError <= io_collectedOutputs_outputs_bits_isError; // @[ReorderBuffer.scala 203:40]
      end else begin
        buffer_12_isError <= _GEN_1390;
      end
    end else begin
      buffer_12_isError <= _GEN_1390;
    end
    if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'hd == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_13_destinationRegister <= io_decoders_0_destination_destinationRegister; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      buffer_13_valueReady <= _GEN_1769;
    end else if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'hd == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_13_valueReady <= 1'h0; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      if (4'hd == io_collectedOutputs_outputs_bits_tag_id) begin // @[ReorderBuffer.scala 202:38]
        buffer_13_value <= io_collectedOutputs_outputs_bits_value; // @[ReorderBuffer.scala 202:38]
      end else begin
        buffer_13_value <= _GEN_1343;
      end
    end else begin
      buffer_13_value <= _GEN_1343;
    end
    if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'hd == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_13_storeSign <= io_decoders_0_destination_storeSign; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      if (4'hd == io_collectedOutputs_outputs_bits_tag_id) begin // @[ReorderBuffer.scala 203:40]
        buffer_13_isError <= io_collectedOutputs_outputs_bits_isError; // @[ReorderBuffer.scala 203:40]
      end else begin
        buffer_13_isError <= _GEN_1391;
      end
    end else begin
      buffer_13_isError <= _GEN_1391;
    end
    if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'he == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_14_destinationRegister <= io_decoders_0_destination_destinationRegister; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      buffer_14_valueReady <= _GEN_1770;
    end else if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'he == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_14_valueReady <= 1'h0; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      if (4'he == io_collectedOutputs_outputs_bits_tag_id) begin // @[ReorderBuffer.scala 202:38]
        buffer_14_value <= io_collectedOutputs_outputs_bits_value; // @[ReorderBuffer.scala 202:38]
      end else begin
        buffer_14_value <= _GEN_1344;
      end
    end else begin
      buffer_14_value <= _GEN_1344;
    end
    if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'he == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_14_storeSign <= io_decoders_0_destination_storeSign; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      if (4'he == io_collectedOutputs_outputs_bits_tag_id) begin // @[ReorderBuffer.scala 203:40]
        buffer_14_isError <= io_collectedOutputs_outputs_bits_isError; // @[ReorderBuffer.scala 203:40]
      end else begin
        buffer_14_isError <= _GEN_1392;
      end
    end else begin
      buffer_14_isError <= _GEN_1392;
    end
    if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'hf == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_15_destinationRegister <= io_decoders_0_destination_destinationRegister; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      buffer_15_valueReady <= _GEN_1771;
    end else if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'hf == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_15_valueReady <= 1'h0; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      if (4'hf == io_collectedOutputs_outputs_bits_tag_id) begin // @[ReorderBuffer.scala 202:38]
        buffer_15_value <= io_collectedOutputs_outputs_bits_value; // @[ReorderBuffer.scala 202:38]
      end else begin
        buffer_15_value <= _GEN_1345;
      end
    end else begin
      buffer_15_value <= _GEN_1345;
    end
    if (io_decoders_0_valid & io_decoders_0_ready) begin // @[ReorderBuffer.scala 130:42]
      if (4'hf == head) begin // @[ReorderBuffer.scala 133:27]
        buffer_15_storeSign <= io_decoders_0_destination_storeSign; // @[ReorderBuffer.scala 133:27]
      end
    end
    if (_T_19) begin // @[ReorderBuffer.scala 201:5]
      if (4'hf == io_collectedOutputs_outputs_bits_tag_id) begin // @[ReorderBuffer.scala 203:40]
        buffer_15_isError <= io_collectedOutputs_outputs_bits_isError; // @[ReorderBuffer.scala 203:40]
      end else begin
        buffer_15_isError <= _GEN_1393;
      end
    end else begin
      buffer_15_isError <= _GEN_1393;
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_1_valid <= 1'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      registerTagMap_1_valid <= _GEN_1395;
    end else if (canCommit_3) begin // @[ReorderBuffer.scala 88:21]
      if (_io_registerFile_3_valid_T) begin // @[ReorderBuffer.scala 89:22]
        registerTagMap_1_valid <= _GEN_1078;
      end else begin
        registerTagMap_1_valid <= _GEN_848;
      end
    end else begin
      registerTagMap_1_valid <= _GEN_848;
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_1_tagId <= 4'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      if (5'h1 == io_decoders_0_destination_destinationRegister) begin // @[ReorderBuffer.scala 149:15]
        registerTagMap_1_tagId <= head; // @[ReorderBuffer.scala 149:15]
      end
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_2_valid <= 1'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      registerTagMap_2_valid <= _GEN_1396;
    end else if (canCommit_3) begin // @[ReorderBuffer.scala 88:21]
      if (_io_registerFile_3_valid_T) begin // @[ReorderBuffer.scala 89:22]
        registerTagMap_2_valid <= _GEN_1079;
      end else begin
        registerTagMap_2_valid <= _GEN_849;
      end
    end else begin
      registerTagMap_2_valid <= _GEN_849;
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_2_tagId <= 4'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      if (5'h2 == io_decoders_0_destination_destinationRegister) begin // @[ReorderBuffer.scala 149:15]
        registerTagMap_2_tagId <= head; // @[ReorderBuffer.scala 149:15]
      end
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_3_valid <= 1'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      registerTagMap_3_valid <= _GEN_1397;
    end else if (canCommit_3) begin // @[ReorderBuffer.scala 88:21]
      if (_io_registerFile_3_valid_T) begin // @[ReorderBuffer.scala 89:22]
        registerTagMap_3_valid <= _GEN_1080;
      end else begin
        registerTagMap_3_valid <= _GEN_850;
      end
    end else begin
      registerTagMap_3_valid <= _GEN_850;
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_3_tagId <= 4'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      if (5'h3 == io_decoders_0_destination_destinationRegister) begin // @[ReorderBuffer.scala 149:15]
        registerTagMap_3_tagId <= head; // @[ReorderBuffer.scala 149:15]
      end
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_4_valid <= 1'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      registerTagMap_4_valid <= _GEN_1398;
    end else if (canCommit_3) begin // @[ReorderBuffer.scala 88:21]
      if (_io_registerFile_3_valid_T) begin // @[ReorderBuffer.scala 89:22]
        registerTagMap_4_valid <= _GEN_1081;
      end else begin
        registerTagMap_4_valid <= _GEN_851;
      end
    end else begin
      registerTagMap_4_valid <= _GEN_851;
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_4_tagId <= 4'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      if (5'h4 == io_decoders_0_destination_destinationRegister) begin // @[ReorderBuffer.scala 149:15]
        registerTagMap_4_tagId <= head; // @[ReorderBuffer.scala 149:15]
      end
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_5_valid <= 1'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      registerTagMap_5_valid <= _GEN_1399;
    end else if (canCommit_3) begin // @[ReorderBuffer.scala 88:21]
      if (_io_registerFile_3_valid_T) begin // @[ReorderBuffer.scala 89:22]
        registerTagMap_5_valid <= _GEN_1082;
      end else begin
        registerTagMap_5_valid <= _GEN_852;
      end
    end else begin
      registerTagMap_5_valid <= _GEN_852;
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_5_tagId <= 4'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      if (5'h5 == io_decoders_0_destination_destinationRegister) begin // @[ReorderBuffer.scala 149:15]
        registerTagMap_5_tagId <= head; // @[ReorderBuffer.scala 149:15]
      end
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_6_valid <= 1'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      registerTagMap_6_valid <= _GEN_1400;
    end else if (canCommit_3) begin // @[ReorderBuffer.scala 88:21]
      if (_io_registerFile_3_valid_T) begin // @[ReorderBuffer.scala 89:22]
        registerTagMap_6_valid <= _GEN_1083;
      end else begin
        registerTagMap_6_valid <= _GEN_853;
      end
    end else begin
      registerTagMap_6_valid <= _GEN_853;
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_6_tagId <= 4'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      if (5'h6 == io_decoders_0_destination_destinationRegister) begin // @[ReorderBuffer.scala 149:15]
        registerTagMap_6_tagId <= head; // @[ReorderBuffer.scala 149:15]
      end
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_7_valid <= 1'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      registerTagMap_7_valid <= _GEN_1401;
    end else if (canCommit_3) begin // @[ReorderBuffer.scala 88:21]
      if (_io_registerFile_3_valid_T) begin // @[ReorderBuffer.scala 89:22]
        registerTagMap_7_valid <= _GEN_1084;
      end else begin
        registerTagMap_7_valid <= _GEN_854;
      end
    end else begin
      registerTagMap_7_valid <= _GEN_854;
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_7_tagId <= 4'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      if (5'h7 == io_decoders_0_destination_destinationRegister) begin // @[ReorderBuffer.scala 149:15]
        registerTagMap_7_tagId <= head; // @[ReorderBuffer.scala 149:15]
      end
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_8_valid <= 1'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      registerTagMap_8_valid <= _GEN_1402;
    end else if (canCommit_3) begin // @[ReorderBuffer.scala 88:21]
      if (_io_registerFile_3_valid_T) begin // @[ReorderBuffer.scala 89:22]
        registerTagMap_8_valid <= _GEN_1085;
      end else begin
        registerTagMap_8_valid <= _GEN_855;
      end
    end else begin
      registerTagMap_8_valid <= _GEN_855;
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_8_tagId <= 4'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      if (5'h8 == io_decoders_0_destination_destinationRegister) begin // @[ReorderBuffer.scala 149:15]
        registerTagMap_8_tagId <= head; // @[ReorderBuffer.scala 149:15]
      end
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_9_valid <= 1'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      registerTagMap_9_valid <= _GEN_1403;
    end else if (canCommit_3) begin // @[ReorderBuffer.scala 88:21]
      if (_io_registerFile_3_valid_T) begin // @[ReorderBuffer.scala 89:22]
        registerTagMap_9_valid <= _GEN_1086;
      end else begin
        registerTagMap_9_valid <= _GEN_856;
      end
    end else begin
      registerTagMap_9_valid <= _GEN_856;
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_9_tagId <= 4'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      if (5'h9 == io_decoders_0_destination_destinationRegister) begin // @[ReorderBuffer.scala 149:15]
        registerTagMap_9_tagId <= head; // @[ReorderBuffer.scala 149:15]
      end
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_10_valid <= 1'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      registerTagMap_10_valid <= _GEN_1404;
    end else if (canCommit_3) begin // @[ReorderBuffer.scala 88:21]
      if (_io_registerFile_3_valid_T) begin // @[ReorderBuffer.scala 89:22]
        registerTagMap_10_valid <= _GEN_1087;
      end else begin
        registerTagMap_10_valid <= _GEN_857;
      end
    end else begin
      registerTagMap_10_valid <= _GEN_857;
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_10_tagId <= 4'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      if (5'ha == io_decoders_0_destination_destinationRegister) begin // @[ReorderBuffer.scala 149:15]
        registerTagMap_10_tagId <= head; // @[ReorderBuffer.scala 149:15]
      end
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_11_valid <= 1'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      registerTagMap_11_valid <= _GEN_1405;
    end else if (canCommit_3) begin // @[ReorderBuffer.scala 88:21]
      if (_io_registerFile_3_valid_T) begin // @[ReorderBuffer.scala 89:22]
        registerTagMap_11_valid <= _GEN_1088;
      end else begin
        registerTagMap_11_valid <= _GEN_858;
      end
    end else begin
      registerTagMap_11_valid <= _GEN_858;
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_11_tagId <= 4'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      if (5'hb == io_decoders_0_destination_destinationRegister) begin // @[ReorderBuffer.scala 149:15]
        registerTagMap_11_tagId <= head; // @[ReorderBuffer.scala 149:15]
      end
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_12_valid <= 1'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      registerTagMap_12_valid <= _GEN_1406;
    end else if (canCommit_3) begin // @[ReorderBuffer.scala 88:21]
      if (_io_registerFile_3_valid_T) begin // @[ReorderBuffer.scala 89:22]
        registerTagMap_12_valid <= _GEN_1089;
      end else begin
        registerTagMap_12_valid <= _GEN_859;
      end
    end else begin
      registerTagMap_12_valid <= _GEN_859;
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_12_tagId <= 4'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      if (5'hc == io_decoders_0_destination_destinationRegister) begin // @[ReorderBuffer.scala 149:15]
        registerTagMap_12_tagId <= head; // @[ReorderBuffer.scala 149:15]
      end
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_13_valid <= 1'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      registerTagMap_13_valid <= _GEN_1407;
    end else if (canCommit_3) begin // @[ReorderBuffer.scala 88:21]
      if (_io_registerFile_3_valid_T) begin // @[ReorderBuffer.scala 89:22]
        registerTagMap_13_valid <= _GEN_1090;
      end else begin
        registerTagMap_13_valid <= _GEN_860;
      end
    end else begin
      registerTagMap_13_valid <= _GEN_860;
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_13_tagId <= 4'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      if (5'hd == io_decoders_0_destination_destinationRegister) begin // @[ReorderBuffer.scala 149:15]
        registerTagMap_13_tagId <= head; // @[ReorderBuffer.scala 149:15]
      end
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_14_valid <= 1'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      registerTagMap_14_valid <= _GEN_1408;
    end else if (canCommit_3) begin // @[ReorderBuffer.scala 88:21]
      if (_io_registerFile_3_valid_T) begin // @[ReorderBuffer.scala 89:22]
        registerTagMap_14_valid <= _GEN_1091;
      end else begin
        registerTagMap_14_valid <= _GEN_861;
      end
    end else begin
      registerTagMap_14_valid <= _GEN_861;
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_14_tagId <= 4'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      if (5'he == io_decoders_0_destination_destinationRegister) begin // @[ReorderBuffer.scala 149:15]
        registerTagMap_14_tagId <= head; // @[ReorderBuffer.scala 149:15]
      end
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_15_valid <= 1'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      registerTagMap_15_valid <= _GEN_1409;
    end else if (canCommit_3) begin // @[ReorderBuffer.scala 88:21]
      if (_io_registerFile_3_valid_T) begin // @[ReorderBuffer.scala 89:22]
        registerTagMap_15_valid <= _GEN_1092;
      end else begin
        registerTagMap_15_valid <= _GEN_862;
      end
    end else begin
      registerTagMap_15_valid <= _GEN_862;
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_15_tagId <= 4'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      if (5'hf == io_decoders_0_destination_destinationRegister) begin // @[ReorderBuffer.scala 149:15]
        registerTagMap_15_tagId <= head; // @[ReorderBuffer.scala 149:15]
      end
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_16_valid <= 1'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      registerTagMap_16_valid <= _GEN_1410;
    end else if (canCommit_3) begin // @[ReorderBuffer.scala 88:21]
      if (_io_registerFile_3_valid_T) begin // @[ReorderBuffer.scala 89:22]
        registerTagMap_16_valid <= _GEN_1093;
      end else begin
        registerTagMap_16_valid <= _GEN_863;
      end
    end else begin
      registerTagMap_16_valid <= _GEN_863;
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_16_tagId <= 4'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      if (5'h10 == io_decoders_0_destination_destinationRegister) begin // @[ReorderBuffer.scala 149:15]
        registerTagMap_16_tagId <= head; // @[ReorderBuffer.scala 149:15]
      end
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_17_valid <= 1'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      registerTagMap_17_valid <= _GEN_1411;
    end else if (canCommit_3) begin // @[ReorderBuffer.scala 88:21]
      if (_io_registerFile_3_valid_T) begin // @[ReorderBuffer.scala 89:22]
        registerTagMap_17_valid <= _GEN_1094;
      end else begin
        registerTagMap_17_valid <= _GEN_864;
      end
    end else begin
      registerTagMap_17_valid <= _GEN_864;
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_17_tagId <= 4'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      if (5'h11 == io_decoders_0_destination_destinationRegister) begin // @[ReorderBuffer.scala 149:15]
        registerTagMap_17_tagId <= head; // @[ReorderBuffer.scala 149:15]
      end
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_18_valid <= 1'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      registerTagMap_18_valid <= _GEN_1412;
    end else if (canCommit_3) begin // @[ReorderBuffer.scala 88:21]
      if (_io_registerFile_3_valid_T) begin // @[ReorderBuffer.scala 89:22]
        registerTagMap_18_valid <= _GEN_1095;
      end else begin
        registerTagMap_18_valid <= _GEN_865;
      end
    end else begin
      registerTagMap_18_valid <= _GEN_865;
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_18_tagId <= 4'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      if (5'h12 == io_decoders_0_destination_destinationRegister) begin // @[ReorderBuffer.scala 149:15]
        registerTagMap_18_tagId <= head; // @[ReorderBuffer.scala 149:15]
      end
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_19_valid <= 1'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      registerTagMap_19_valid <= _GEN_1413;
    end else if (canCommit_3) begin // @[ReorderBuffer.scala 88:21]
      if (_io_registerFile_3_valid_T) begin // @[ReorderBuffer.scala 89:22]
        registerTagMap_19_valid <= _GEN_1096;
      end else begin
        registerTagMap_19_valid <= _GEN_866;
      end
    end else begin
      registerTagMap_19_valid <= _GEN_866;
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_19_tagId <= 4'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      if (5'h13 == io_decoders_0_destination_destinationRegister) begin // @[ReorderBuffer.scala 149:15]
        registerTagMap_19_tagId <= head; // @[ReorderBuffer.scala 149:15]
      end
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_20_valid <= 1'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      registerTagMap_20_valid <= _GEN_1414;
    end else if (canCommit_3) begin // @[ReorderBuffer.scala 88:21]
      if (_io_registerFile_3_valid_T) begin // @[ReorderBuffer.scala 89:22]
        registerTagMap_20_valid <= _GEN_1097;
      end else begin
        registerTagMap_20_valid <= _GEN_867;
      end
    end else begin
      registerTagMap_20_valid <= _GEN_867;
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_20_tagId <= 4'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      if (5'h14 == io_decoders_0_destination_destinationRegister) begin // @[ReorderBuffer.scala 149:15]
        registerTagMap_20_tagId <= head; // @[ReorderBuffer.scala 149:15]
      end
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_21_valid <= 1'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      registerTagMap_21_valid <= _GEN_1415;
    end else if (canCommit_3) begin // @[ReorderBuffer.scala 88:21]
      if (_io_registerFile_3_valid_T) begin // @[ReorderBuffer.scala 89:22]
        registerTagMap_21_valid <= _GEN_1098;
      end else begin
        registerTagMap_21_valid <= _GEN_868;
      end
    end else begin
      registerTagMap_21_valid <= _GEN_868;
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_21_tagId <= 4'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      if (5'h15 == io_decoders_0_destination_destinationRegister) begin // @[ReorderBuffer.scala 149:15]
        registerTagMap_21_tagId <= head; // @[ReorderBuffer.scala 149:15]
      end
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_22_valid <= 1'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      registerTagMap_22_valid <= _GEN_1416;
    end else if (canCommit_3) begin // @[ReorderBuffer.scala 88:21]
      if (_io_registerFile_3_valid_T) begin // @[ReorderBuffer.scala 89:22]
        registerTagMap_22_valid <= _GEN_1099;
      end else begin
        registerTagMap_22_valid <= _GEN_869;
      end
    end else begin
      registerTagMap_22_valid <= _GEN_869;
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_22_tagId <= 4'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      if (5'h16 == io_decoders_0_destination_destinationRegister) begin // @[ReorderBuffer.scala 149:15]
        registerTagMap_22_tagId <= head; // @[ReorderBuffer.scala 149:15]
      end
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_23_valid <= 1'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      registerTagMap_23_valid <= _GEN_1417;
    end else if (canCommit_3) begin // @[ReorderBuffer.scala 88:21]
      if (_io_registerFile_3_valid_T) begin // @[ReorderBuffer.scala 89:22]
        registerTagMap_23_valid <= _GEN_1100;
      end else begin
        registerTagMap_23_valid <= _GEN_870;
      end
    end else begin
      registerTagMap_23_valid <= _GEN_870;
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_23_tagId <= 4'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      if (5'h17 == io_decoders_0_destination_destinationRegister) begin // @[ReorderBuffer.scala 149:15]
        registerTagMap_23_tagId <= head; // @[ReorderBuffer.scala 149:15]
      end
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_24_valid <= 1'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      registerTagMap_24_valid <= _GEN_1418;
    end else if (canCommit_3) begin // @[ReorderBuffer.scala 88:21]
      if (_io_registerFile_3_valid_T) begin // @[ReorderBuffer.scala 89:22]
        registerTagMap_24_valid <= _GEN_1101;
      end else begin
        registerTagMap_24_valid <= _GEN_871;
      end
    end else begin
      registerTagMap_24_valid <= _GEN_871;
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_24_tagId <= 4'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      if (5'h18 == io_decoders_0_destination_destinationRegister) begin // @[ReorderBuffer.scala 149:15]
        registerTagMap_24_tagId <= head; // @[ReorderBuffer.scala 149:15]
      end
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_25_valid <= 1'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      registerTagMap_25_valid <= _GEN_1419;
    end else if (canCommit_3) begin // @[ReorderBuffer.scala 88:21]
      if (_io_registerFile_3_valid_T) begin // @[ReorderBuffer.scala 89:22]
        registerTagMap_25_valid <= _GEN_1102;
      end else begin
        registerTagMap_25_valid <= _GEN_872;
      end
    end else begin
      registerTagMap_25_valid <= _GEN_872;
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_25_tagId <= 4'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      if (5'h19 == io_decoders_0_destination_destinationRegister) begin // @[ReorderBuffer.scala 149:15]
        registerTagMap_25_tagId <= head; // @[ReorderBuffer.scala 149:15]
      end
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_26_valid <= 1'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      registerTagMap_26_valid <= _GEN_1420;
    end else if (canCommit_3) begin // @[ReorderBuffer.scala 88:21]
      if (_io_registerFile_3_valid_T) begin // @[ReorderBuffer.scala 89:22]
        registerTagMap_26_valid <= _GEN_1103;
      end else begin
        registerTagMap_26_valid <= _GEN_873;
      end
    end else begin
      registerTagMap_26_valid <= _GEN_873;
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_26_tagId <= 4'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      if (5'h1a == io_decoders_0_destination_destinationRegister) begin // @[ReorderBuffer.scala 149:15]
        registerTagMap_26_tagId <= head; // @[ReorderBuffer.scala 149:15]
      end
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_27_valid <= 1'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      registerTagMap_27_valid <= _GEN_1421;
    end else if (canCommit_3) begin // @[ReorderBuffer.scala 88:21]
      if (_io_registerFile_3_valid_T) begin // @[ReorderBuffer.scala 89:22]
        registerTagMap_27_valid <= _GEN_1104;
      end else begin
        registerTagMap_27_valid <= _GEN_874;
      end
    end else begin
      registerTagMap_27_valid <= _GEN_874;
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_27_tagId <= 4'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      if (5'h1b == io_decoders_0_destination_destinationRegister) begin // @[ReorderBuffer.scala 149:15]
        registerTagMap_27_tagId <= head; // @[ReorderBuffer.scala 149:15]
      end
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_28_valid <= 1'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      registerTagMap_28_valid <= _GEN_1422;
    end else if (canCommit_3) begin // @[ReorderBuffer.scala 88:21]
      if (_io_registerFile_3_valid_T) begin // @[ReorderBuffer.scala 89:22]
        registerTagMap_28_valid <= _GEN_1105;
      end else begin
        registerTagMap_28_valid <= _GEN_875;
      end
    end else begin
      registerTagMap_28_valid <= _GEN_875;
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_28_tagId <= 4'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      if (5'h1c == io_decoders_0_destination_destinationRegister) begin // @[ReorderBuffer.scala 149:15]
        registerTagMap_28_tagId <= head; // @[ReorderBuffer.scala 149:15]
      end
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_29_valid <= 1'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      registerTagMap_29_valid <= _GEN_1423;
    end else if (canCommit_3) begin // @[ReorderBuffer.scala 88:21]
      if (_io_registerFile_3_valid_T) begin // @[ReorderBuffer.scala 89:22]
        registerTagMap_29_valid <= _GEN_1106;
      end else begin
        registerTagMap_29_valid <= _GEN_876;
      end
    end else begin
      registerTagMap_29_valid <= _GEN_876;
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_29_tagId <= 4'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      if (5'h1d == io_decoders_0_destination_destinationRegister) begin // @[ReorderBuffer.scala 149:15]
        registerTagMap_29_tagId <= head; // @[ReorderBuffer.scala 149:15]
      end
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_30_valid <= 1'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      registerTagMap_30_valid <= _GEN_1424;
    end else if (canCommit_3) begin // @[ReorderBuffer.scala 88:21]
      if (_io_registerFile_3_valid_T) begin // @[ReorderBuffer.scala 89:22]
        registerTagMap_30_valid <= _GEN_1107;
      end else begin
        registerTagMap_30_valid <= _GEN_877;
      end
    end else begin
      registerTagMap_30_valid <= _GEN_877;
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_30_tagId <= 4'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      if (5'h1e == io_decoders_0_destination_destinationRegister) begin // @[ReorderBuffer.scala 149:15]
        registerTagMap_30_tagId <= head; // @[ReorderBuffer.scala 149:15]
      end
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_31_valid <= 1'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      registerTagMap_31_valid <= _GEN_1425;
    end else if (canCommit_3) begin // @[ReorderBuffer.scala 88:21]
      if (_io_registerFile_3_valid_T) begin // @[ReorderBuffer.scala 89:22]
        registerTagMap_31_valid <= _GEN_1108;
      end else begin
        registerTagMap_31_valid <= _GEN_878;
      end
    end else begin
      registerTagMap_31_valid <= _GEN_878;
    end
    if (reset) begin // @[ReorderBuffer.scala 69:39]
      registerTagMap_31_tagId <= 4'h0; // @[ReorderBuffer.scala 69:39]
    end else if (io_decoders_0_destination_destinationRegister != 5'h0) begin // @[ReorderBuffer.scala 145:59]
      if (5'h1f == io_decoders_0_destination_destinationRegister) begin // @[ReorderBuffer.scala 149:15]
        registerTagMap_31_tagId <= head; // @[ReorderBuffer.scala 149:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  head = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  tail = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  buffer_0_destinationRegister = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  buffer_0_valueReady = _RAND_3[0:0];
  _RAND_4 = {2{`RANDOM}};
  buffer_0_value = _RAND_4[63:0];
  _RAND_5 = {1{`RANDOM}};
  buffer_0_storeSign = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  buffer_0_isError = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  buffer_1_destinationRegister = _RAND_7[4:0];
  _RAND_8 = {1{`RANDOM}};
  buffer_1_valueReady = _RAND_8[0:0];
  _RAND_9 = {2{`RANDOM}};
  buffer_1_value = _RAND_9[63:0];
  _RAND_10 = {1{`RANDOM}};
  buffer_1_storeSign = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  buffer_1_isError = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  buffer_2_destinationRegister = _RAND_12[4:0];
  _RAND_13 = {1{`RANDOM}};
  buffer_2_valueReady = _RAND_13[0:0];
  _RAND_14 = {2{`RANDOM}};
  buffer_2_value = _RAND_14[63:0];
  _RAND_15 = {1{`RANDOM}};
  buffer_2_storeSign = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  buffer_2_isError = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  buffer_3_destinationRegister = _RAND_17[4:0];
  _RAND_18 = {1{`RANDOM}};
  buffer_3_valueReady = _RAND_18[0:0];
  _RAND_19 = {2{`RANDOM}};
  buffer_3_value = _RAND_19[63:0];
  _RAND_20 = {1{`RANDOM}};
  buffer_3_storeSign = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  buffer_3_isError = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  buffer_4_destinationRegister = _RAND_22[4:0];
  _RAND_23 = {1{`RANDOM}};
  buffer_4_valueReady = _RAND_23[0:0];
  _RAND_24 = {2{`RANDOM}};
  buffer_4_value = _RAND_24[63:0];
  _RAND_25 = {1{`RANDOM}};
  buffer_4_storeSign = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  buffer_4_isError = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  buffer_5_destinationRegister = _RAND_27[4:0];
  _RAND_28 = {1{`RANDOM}};
  buffer_5_valueReady = _RAND_28[0:0];
  _RAND_29 = {2{`RANDOM}};
  buffer_5_value = _RAND_29[63:0];
  _RAND_30 = {1{`RANDOM}};
  buffer_5_storeSign = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  buffer_5_isError = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  buffer_6_destinationRegister = _RAND_32[4:0];
  _RAND_33 = {1{`RANDOM}};
  buffer_6_valueReady = _RAND_33[0:0];
  _RAND_34 = {2{`RANDOM}};
  buffer_6_value = _RAND_34[63:0];
  _RAND_35 = {1{`RANDOM}};
  buffer_6_storeSign = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  buffer_6_isError = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  buffer_7_destinationRegister = _RAND_37[4:0];
  _RAND_38 = {1{`RANDOM}};
  buffer_7_valueReady = _RAND_38[0:0];
  _RAND_39 = {2{`RANDOM}};
  buffer_7_value = _RAND_39[63:0];
  _RAND_40 = {1{`RANDOM}};
  buffer_7_storeSign = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  buffer_7_isError = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  buffer_8_destinationRegister = _RAND_42[4:0];
  _RAND_43 = {1{`RANDOM}};
  buffer_8_valueReady = _RAND_43[0:0];
  _RAND_44 = {2{`RANDOM}};
  buffer_8_value = _RAND_44[63:0];
  _RAND_45 = {1{`RANDOM}};
  buffer_8_storeSign = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  buffer_8_isError = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  buffer_9_destinationRegister = _RAND_47[4:0];
  _RAND_48 = {1{`RANDOM}};
  buffer_9_valueReady = _RAND_48[0:0];
  _RAND_49 = {2{`RANDOM}};
  buffer_9_value = _RAND_49[63:0];
  _RAND_50 = {1{`RANDOM}};
  buffer_9_storeSign = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  buffer_9_isError = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  buffer_10_destinationRegister = _RAND_52[4:0];
  _RAND_53 = {1{`RANDOM}};
  buffer_10_valueReady = _RAND_53[0:0];
  _RAND_54 = {2{`RANDOM}};
  buffer_10_value = _RAND_54[63:0];
  _RAND_55 = {1{`RANDOM}};
  buffer_10_storeSign = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  buffer_10_isError = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  buffer_11_destinationRegister = _RAND_57[4:0];
  _RAND_58 = {1{`RANDOM}};
  buffer_11_valueReady = _RAND_58[0:0];
  _RAND_59 = {2{`RANDOM}};
  buffer_11_value = _RAND_59[63:0];
  _RAND_60 = {1{`RANDOM}};
  buffer_11_storeSign = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  buffer_11_isError = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  buffer_12_destinationRegister = _RAND_62[4:0];
  _RAND_63 = {1{`RANDOM}};
  buffer_12_valueReady = _RAND_63[0:0];
  _RAND_64 = {2{`RANDOM}};
  buffer_12_value = _RAND_64[63:0];
  _RAND_65 = {1{`RANDOM}};
  buffer_12_storeSign = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  buffer_12_isError = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  buffer_13_destinationRegister = _RAND_67[4:0];
  _RAND_68 = {1{`RANDOM}};
  buffer_13_valueReady = _RAND_68[0:0];
  _RAND_69 = {2{`RANDOM}};
  buffer_13_value = _RAND_69[63:0];
  _RAND_70 = {1{`RANDOM}};
  buffer_13_storeSign = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  buffer_13_isError = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  buffer_14_destinationRegister = _RAND_72[4:0];
  _RAND_73 = {1{`RANDOM}};
  buffer_14_valueReady = _RAND_73[0:0];
  _RAND_74 = {2{`RANDOM}};
  buffer_14_value = _RAND_74[63:0];
  _RAND_75 = {1{`RANDOM}};
  buffer_14_storeSign = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  buffer_14_isError = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  buffer_15_destinationRegister = _RAND_77[4:0];
  _RAND_78 = {1{`RANDOM}};
  buffer_15_valueReady = _RAND_78[0:0];
  _RAND_79 = {2{`RANDOM}};
  buffer_15_value = _RAND_79[63:0];
  _RAND_80 = {1{`RANDOM}};
  buffer_15_storeSign = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  buffer_15_isError = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  registerTagMap_1_valid = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  registerTagMap_1_tagId = _RAND_83[3:0];
  _RAND_84 = {1{`RANDOM}};
  registerTagMap_2_valid = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  registerTagMap_2_tagId = _RAND_85[3:0];
  _RAND_86 = {1{`RANDOM}};
  registerTagMap_3_valid = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  registerTagMap_3_tagId = _RAND_87[3:0];
  _RAND_88 = {1{`RANDOM}};
  registerTagMap_4_valid = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  registerTagMap_4_tagId = _RAND_89[3:0];
  _RAND_90 = {1{`RANDOM}};
  registerTagMap_5_valid = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  registerTagMap_5_tagId = _RAND_91[3:0];
  _RAND_92 = {1{`RANDOM}};
  registerTagMap_6_valid = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  registerTagMap_6_tagId = _RAND_93[3:0];
  _RAND_94 = {1{`RANDOM}};
  registerTagMap_7_valid = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  registerTagMap_7_tagId = _RAND_95[3:0];
  _RAND_96 = {1{`RANDOM}};
  registerTagMap_8_valid = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  registerTagMap_8_tagId = _RAND_97[3:0];
  _RAND_98 = {1{`RANDOM}};
  registerTagMap_9_valid = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  registerTagMap_9_tagId = _RAND_99[3:0];
  _RAND_100 = {1{`RANDOM}};
  registerTagMap_10_valid = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  registerTagMap_10_tagId = _RAND_101[3:0];
  _RAND_102 = {1{`RANDOM}};
  registerTagMap_11_valid = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  registerTagMap_11_tagId = _RAND_103[3:0];
  _RAND_104 = {1{`RANDOM}};
  registerTagMap_12_valid = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  registerTagMap_12_tagId = _RAND_105[3:0];
  _RAND_106 = {1{`RANDOM}};
  registerTagMap_13_valid = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  registerTagMap_13_tagId = _RAND_107[3:0];
  _RAND_108 = {1{`RANDOM}};
  registerTagMap_14_valid = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  registerTagMap_14_tagId = _RAND_109[3:0];
  _RAND_110 = {1{`RANDOM}};
  registerTagMap_15_valid = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  registerTagMap_15_tagId = _RAND_111[3:0];
  _RAND_112 = {1{`RANDOM}};
  registerTagMap_16_valid = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  registerTagMap_16_tagId = _RAND_113[3:0];
  _RAND_114 = {1{`RANDOM}};
  registerTagMap_17_valid = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  registerTagMap_17_tagId = _RAND_115[3:0];
  _RAND_116 = {1{`RANDOM}};
  registerTagMap_18_valid = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  registerTagMap_18_tagId = _RAND_117[3:0];
  _RAND_118 = {1{`RANDOM}};
  registerTagMap_19_valid = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  registerTagMap_19_tagId = _RAND_119[3:0];
  _RAND_120 = {1{`RANDOM}};
  registerTagMap_20_valid = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  registerTagMap_20_tagId = _RAND_121[3:0];
  _RAND_122 = {1{`RANDOM}};
  registerTagMap_21_valid = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  registerTagMap_21_tagId = _RAND_123[3:0];
  _RAND_124 = {1{`RANDOM}};
  registerTagMap_22_valid = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  registerTagMap_22_tagId = _RAND_125[3:0];
  _RAND_126 = {1{`RANDOM}};
  registerTagMap_23_valid = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  registerTagMap_23_tagId = _RAND_127[3:0];
  _RAND_128 = {1{`RANDOM}};
  registerTagMap_24_valid = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  registerTagMap_24_tagId = _RAND_129[3:0];
  _RAND_130 = {1{`RANDOM}};
  registerTagMap_25_valid = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  registerTagMap_25_tagId = _RAND_131[3:0];
  _RAND_132 = {1{`RANDOM}};
  registerTagMap_26_valid = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  registerTagMap_26_tagId = _RAND_133[3:0];
  _RAND_134 = {1{`RANDOM}};
  registerTagMap_27_valid = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  registerTagMap_27_tagId = _RAND_135[3:0];
  _RAND_136 = {1{`RANDOM}};
  registerTagMap_28_valid = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  registerTagMap_28_tagId = _RAND_137[3:0];
  _RAND_138 = {1{`RANDOM}};
  registerTagMap_29_valid = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  registerTagMap_29_tagId = _RAND_139[3:0];
  _RAND_140 = {1{`RANDOM}};
  registerTagMap_30_valid = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  registerTagMap_30_tagId = _RAND_141[3:0];
  _RAND_142 = {1{`RANDOM}};
  registerTagMap_31_valid = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  registerTagMap_31_tagId = _RAND_143[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RegisterFile(
  input         clock,
  input         reset,
  input  [4:0]  io_decoders_0_sourceRegister1,
  input  [4:0]  io_decoders_0_sourceRegister2,
  output [63:0] io_decoders_0_value1,
  output [63:0] io_decoders_0_value2,
  input         io_reorderBuffer_0_valid,
  input  [4:0]  io_reorderBuffer_0_bits_destinationRegister,
  input  [63:0] io_reorderBuffer_0_bits_value,
  input         io_reorderBuffer_1_valid,
  input  [4:0]  io_reorderBuffer_1_bits_destinationRegister,
  input  [63:0] io_reorderBuffer_1_bits_value,
  input         io_reorderBuffer_2_valid,
  input  [4:0]  io_reorderBuffer_2_bits_destinationRegister,
  input  [63:0] io_reorderBuffer_2_bits_value,
  input         io_reorderBuffer_3_valid,
  input  [4:0]  io_reorderBuffer_3_bits_destinationRegister,
  input  [63:0] io_reorderBuffer_3_bits_value
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] registers_1; // @[RegisterFile.scala 37:26]
  reg [63:0] registers_2; // @[RegisterFile.scala 37:26]
  reg [63:0] registers_3; // @[RegisterFile.scala 37:26]
  reg [63:0] registers_4; // @[RegisterFile.scala 37:26]
  reg [63:0] registers_5; // @[RegisterFile.scala 37:26]
  reg [63:0] registers_6; // @[RegisterFile.scala 37:26]
  reg [63:0] registers_7; // @[RegisterFile.scala 37:26]
  reg [63:0] registers_8; // @[RegisterFile.scala 37:26]
  reg [63:0] registers_9; // @[RegisterFile.scala 37:26]
  reg [63:0] registers_10; // @[RegisterFile.scala 37:26]
  reg [63:0] registers_11; // @[RegisterFile.scala 37:26]
  reg [63:0] registers_12; // @[RegisterFile.scala 37:26]
  reg [63:0] registers_13; // @[RegisterFile.scala 37:26]
  reg [63:0] registers_14; // @[RegisterFile.scala 37:26]
  reg [63:0] registers_15; // @[RegisterFile.scala 37:26]
  reg [63:0] registers_16; // @[RegisterFile.scala 37:26]
  reg [63:0] registers_17; // @[RegisterFile.scala 37:26]
  reg [63:0] registers_18; // @[RegisterFile.scala 37:26]
  reg [63:0] registers_19; // @[RegisterFile.scala 37:26]
  reg [63:0] registers_20; // @[RegisterFile.scala 37:26]
  reg [63:0] registers_21; // @[RegisterFile.scala 37:26]
  reg [63:0] registers_22; // @[RegisterFile.scala 37:26]
  reg [63:0] registers_23; // @[RegisterFile.scala 37:26]
  reg [63:0] registers_24; // @[RegisterFile.scala 37:26]
  reg [63:0] registers_25; // @[RegisterFile.scala 37:26]
  reg [63:0] registers_26; // @[RegisterFile.scala 37:26]
  reg [63:0] registers_27; // @[RegisterFile.scala 37:26]
  reg [63:0] registers_28; // @[RegisterFile.scala 37:26]
  reg [63:0] registers_29; // @[RegisterFile.scala 37:26]
  reg [63:0] registers_30; // @[RegisterFile.scala 37:26]
  reg [63:0] registers_31; // @[RegisterFile.scala 37:26]
  wire [63:0] _GEN_1 = 5'h1 == io_reorderBuffer_0_bits_destinationRegister ? io_reorderBuffer_0_bits_value : registers_1
    ; // @[RegisterFile.scala 37:26 46:{46,46}]
  wire [63:0] _GEN_2 = 5'h2 == io_reorderBuffer_0_bits_destinationRegister ? io_reorderBuffer_0_bits_value : registers_2
    ; // @[RegisterFile.scala 37:26 46:{46,46}]
  wire [63:0] _GEN_3 = 5'h3 == io_reorderBuffer_0_bits_destinationRegister ? io_reorderBuffer_0_bits_value : registers_3
    ; // @[RegisterFile.scala 37:26 46:{46,46}]
  wire [63:0] _GEN_4 = 5'h4 == io_reorderBuffer_0_bits_destinationRegister ? io_reorderBuffer_0_bits_value : registers_4
    ; // @[RegisterFile.scala 37:26 46:{46,46}]
  wire [63:0] _GEN_5 = 5'h5 == io_reorderBuffer_0_bits_destinationRegister ? io_reorderBuffer_0_bits_value : registers_5
    ; // @[RegisterFile.scala 37:26 46:{46,46}]
  wire [63:0] _GEN_6 = 5'h6 == io_reorderBuffer_0_bits_destinationRegister ? io_reorderBuffer_0_bits_value : registers_6
    ; // @[RegisterFile.scala 37:26 46:{46,46}]
  wire [63:0] _GEN_7 = 5'h7 == io_reorderBuffer_0_bits_destinationRegister ? io_reorderBuffer_0_bits_value : registers_7
    ; // @[RegisterFile.scala 37:26 46:{46,46}]
  wire [63:0] _GEN_8 = 5'h8 == io_reorderBuffer_0_bits_destinationRegister ? io_reorderBuffer_0_bits_value : registers_8
    ; // @[RegisterFile.scala 37:26 46:{46,46}]
  wire [63:0] _GEN_9 = 5'h9 == io_reorderBuffer_0_bits_destinationRegister ? io_reorderBuffer_0_bits_value : registers_9
    ; // @[RegisterFile.scala 37:26 46:{46,46}]
  wire [63:0] _GEN_10 = 5'ha == io_reorderBuffer_0_bits_destinationRegister ? io_reorderBuffer_0_bits_value :
    registers_10; // @[RegisterFile.scala 37:26 46:{46,46}]
  wire [63:0] _GEN_11 = 5'hb == io_reorderBuffer_0_bits_destinationRegister ? io_reorderBuffer_0_bits_value :
    registers_11; // @[RegisterFile.scala 37:26 46:{46,46}]
  wire [63:0] _GEN_12 = 5'hc == io_reorderBuffer_0_bits_destinationRegister ? io_reorderBuffer_0_bits_value :
    registers_12; // @[RegisterFile.scala 37:26 46:{46,46}]
  wire [63:0] _GEN_13 = 5'hd == io_reorderBuffer_0_bits_destinationRegister ? io_reorderBuffer_0_bits_value :
    registers_13; // @[RegisterFile.scala 37:26 46:{46,46}]
  wire [63:0] _GEN_14 = 5'he == io_reorderBuffer_0_bits_destinationRegister ? io_reorderBuffer_0_bits_value :
    registers_14; // @[RegisterFile.scala 37:26 46:{46,46}]
  wire [63:0] _GEN_15 = 5'hf == io_reorderBuffer_0_bits_destinationRegister ? io_reorderBuffer_0_bits_value :
    registers_15; // @[RegisterFile.scala 37:26 46:{46,46}]
  wire [63:0] _GEN_16 = 5'h10 == io_reorderBuffer_0_bits_destinationRegister ? io_reorderBuffer_0_bits_value :
    registers_16; // @[RegisterFile.scala 37:26 46:{46,46}]
  wire [63:0] _GEN_17 = 5'h11 == io_reorderBuffer_0_bits_destinationRegister ? io_reorderBuffer_0_bits_value :
    registers_17; // @[RegisterFile.scala 37:26 46:{46,46}]
  wire [63:0] _GEN_18 = 5'h12 == io_reorderBuffer_0_bits_destinationRegister ? io_reorderBuffer_0_bits_value :
    registers_18; // @[RegisterFile.scala 37:26 46:{46,46}]
  wire [63:0] _GEN_19 = 5'h13 == io_reorderBuffer_0_bits_destinationRegister ? io_reorderBuffer_0_bits_value :
    registers_19; // @[RegisterFile.scala 37:26 46:{46,46}]
  wire [63:0] _GEN_20 = 5'h14 == io_reorderBuffer_0_bits_destinationRegister ? io_reorderBuffer_0_bits_value :
    registers_20; // @[RegisterFile.scala 37:26 46:{46,46}]
  wire [63:0] _GEN_21 = 5'h15 == io_reorderBuffer_0_bits_destinationRegister ? io_reorderBuffer_0_bits_value :
    registers_21; // @[RegisterFile.scala 37:26 46:{46,46}]
  wire [63:0] _GEN_22 = 5'h16 == io_reorderBuffer_0_bits_destinationRegister ? io_reorderBuffer_0_bits_value :
    registers_22; // @[RegisterFile.scala 37:26 46:{46,46}]
  wire [63:0] _GEN_23 = 5'h17 == io_reorderBuffer_0_bits_destinationRegister ? io_reorderBuffer_0_bits_value :
    registers_23; // @[RegisterFile.scala 37:26 46:{46,46}]
  wire [63:0] _GEN_24 = 5'h18 == io_reorderBuffer_0_bits_destinationRegister ? io_reorderBuffer_0_bits_value :
    registers_24; // @[RegisterFile.scala 37:26 46:{46,46}]
  wire [63:0] _GEN_25 = 5'h19 == io_reorderBuffer_0_bits_destinationRegister ? io_reorderBuffer_0_bits_value :
    registers_25; // @[RegisterFile.scala 37:26 46:{46,46}]
  wire [63:0] _GEN_26 = 5'h1a == io_reorderBuffer_0_bits_destinationRegister ? io_reorderBuffer_0_bits_value :
    registers_26; // @[RegisterFile.scala 37:26 46:{46,46}]
  wire [63:0] _GEN_27 = 5'h1b == io_reorderBuffer_0_bits_destinationRegister ? io_reorderBuffer_0_bits_value :
    registers_27; // @[RegisterFile.scala 37:26 46:{46,46}]
  wire [63:0] _GEN_28 = 5'h1c == io_reorderBuffer_0_bits_destinationRegister ? io_reorderBuffer_0_bits_value :
    registers_28; // @[RegisterFile.scala 37:26 46:{46,46}]
  wire [63:0] _GEN_29 = 5'h1d == io_reorderBuffer_0_bits_destinationRegister ? io_reorderBuffer_0_bits_value :
    registers_29; // @[RegisterFile.scala 37:26 46:{46,46}]
  wire [63:0] _GEN_30 = 5'h1e == io_reorderBuffer_0_bits_destinationRegister ? io_reorderBuffer_0_bits_value :
    registers_30; // @[RegisterFile.scala 37:26 46:{46,46}]
  wire [63:0] _GEN_31 = 5'h1f == io_reorderBuffer_0_bits_destinationRegister ? io_reorderBuffer_0_bits_value :
    registers_31; // @[RegisterFile.scala 37:26 46:{46,46}]
  wire [63:0] _GEN_33 = io_reorderBuffer_0_valid ? _GEN_1 : registers_1; // @[RegisterFile.scala 45:20 37:26]
  wire [63:0] _GEN_34 = io_reorderBuffer_0_valid ? _GEN_2 : registers_2; // @[RegisterFile.scala 45:20 37:26]
  wire [63:0] _GEN_35 = io_reorderBuffer_0_valid ? _GEN_3 : registers_3; // @[RegisterFile.scala 45:20 37:26]
  wire [63:0] _GEN_36 = io_reorderBuffer_0_valid ? _GEN_4 : registers_4; // @[RegisterFile.scala 45:20 37:26]
  wire [63:0] _GEN_37 = io_reorderBuffer_0_valid ? _GEN_5 : registers_5; // @[RegisterFile.scala 45:20 37:26]
  wire [63:0] _GEN_38 = io_reorderBuffer_0_valid ? _GEN_6 : registers_6; // @[RegisterFile.scala 45:20 37:26]
  wire [63:0] _GEN_39 = io_reorderBuffer_0_valid ? _GEN_7 : registers_7; // @[RegisterFile.scala 45:20 37:26]
  wire [63:0] _GEN_40 = io_reorderBuffer_0_valid ? _GEN_8 : registers_8; // @[RegisterFile.scala 45:20 37:26]
  wire [63:0] _GEN_41 = io_reorderBuffer_0_valid ? _GEN_9 : registers_9; // @[RegisterFile.scala 45:20 37:26]
  wire [63:0] _GEN_42 = io_reorderBuffer_0_valid ? _GEN_10 : registers_10; // @[RegisterFile.scala 45:20 37:26]
  wire [63:0] _GEN_43 = io_reorderBuffer_0_valid ? _GEN_11 : registers_11; // @[RegisterFile.scala 45:20 37:26]
  wire [63:0] _GEN_44 = io_reorderBuffer_0_valid ? _GEN_12 : registers_12; // @[RegisterFile.scala 45:20 37:26]
  wire [63:0] _GEN_45 = io_reorderBuffer_0_valid ? _GEN_13 : registers_13; // @[RegisterFile.scala 45:20 37:26]
  wire [63:0] _GEN_46 = io_reorderBuffer_0_valid ? _GEN_14 : registers_14; // @[RegisterFile.scala 45:20 37:26]
  wire [63:0] _GEN_47 = io_reorderBuffer_0_valid ? _GEN_15 : registers_15; // @[RegisterFile.scala 45:20 37:26]
  wire [63:0] _GEN_48 = io_reorderBuffer_0_valid ? _GEN_16 : registers_16; // @[RegisterFile.scala 45:20 37:26]
  wire [63:0] _GEN_49 = io_reorderBuffer_0_valid ? _GEN_17 : registers_17; // @[RegisterFile.scala 45:20 37:26]
  wire [63:0] _GEN_50 = io_reorderBuffer_0_valid ? _GEN_18 : registers_18; // @[RegisterFile.scala 45:20 37:26]
  wire [63:0] _GEN_51 = io_reorderBuffer_0_valid ? _GEN_19 : registers_19; // @[RegisterFile.scala 45:20 37:26]
  wire [63:0] _GEN_52 = io_reorderBuffer_0_valid ? _GEN_20 : registers_20; // @[RegisterFile.scala 45:20 37:26]
  wire [63:0] _GEN_53 = io_reorderBuffer_0_valid ? _GEN_21 : registers_21; // @[RegisterFile.scala 45:20 37:26]
  wire [63:0] _GEN_54 = io_reorderBuffer_0_valid ? _GEN_22 : registers_22; // @[RegisterFile.scala 45:20 37:26]
  wire [63:0] _GEN_55 = io_reorderBuffer_0_valid ? _GEN_23 : registers_23; // @[RegisterFile.scala 45:20 37:26]
  wire [63:0] _GEN_56 = io_reorderBuffer_0_valid ? _GEN_24 : registers_24; // @[RegisterFile.scala 45:20 37:26]
  wire [63:0] _GEN_57 = io_reorderBuffer_0_valid ? _GEN_25 : registers_25; // @[RegisterFile.scala 45:20 37:26]
  wire [63:0] _GEN_58 = io_reorderBuffer_0_valid ? _GEN_26 : registers_26; // @[RegisterFile.scala 45:20 37:26]
  wire [63:0] _GEN_59 = io_reorderBuffer_0_valid ? _GEN_27 : registers_27; // @[RegisterFile.scala 45:20 37:26]
  wire [63:0] _GEN_60 = io_reorderBuffer_0_valid ? _GEN_28 : registers_28; // @[RegisterFile.scala 45:20 37:26]
  wire [63:0] _GEN_61 = io_reorderBuffer_0_valid ? _GEN_29 : registers_29; // @[RegisterFile.scala 45:20 37:26]
  wire [63:0] _GEN_62 = io_reorderBuffer_0_valid ? _GEN_30 : registers_30; // @[RegisterFile.scala 45:20 37:26]
  wire [63:0] _GEN_63 = io_reorderBuffer_0_valid ? _GEN_31 : registers_31; // @[RegisterFile.scala 45:20 37:26]
  wire [63:0] _GEN_65 = 5'h1 == io_reorderBuffer_1_bits_destinationRegister ? io_reorderBuffer_1_bits_value : _GEN_33; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_66 = 5'h2 == io_reorderBuffer_1_bits_destinationRegister ? io_reorderBuffer_1_bits_value : _GEN_34; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_67 = 5'h3 == io_reorderBuffer_1_bits_destinationRegister ? io_reorderBuffer_1_bits_value : _GEN_35; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_68 = 5'h4 == io_reorderBuffer_1_bits_destinationRegister ? io_reorderBuffer_1_bits_value : _GEN_36; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_69 = 5'h5 == io_reorderBuffer_1_bits_destinationRegister ? io_reorderBuffer_1_bits_value : _GEN_37; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_70 = 5'h6 == io_reorderBuffer_1_bits_destinationRegister ? io_reorderBuffer_1_bits_value : _GEN_38; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_71 = 5'h7 == io_reorderBuffer_1_bits_destinationRegister ? io_reorderBuffer_1_bits_value : _GEN_39; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_72 = 5'h8 == io_reorderBuffer_1_bits_destinationRegister ? io_reorderBuffer_1_bits_value : _GEN_40; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_73 = 5'h9 == io_reorderBuffer_1_bits_destinationRegister ? io_reorderBuffer_1_bits_value : _GEN_41; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_74 = 5'ha == io_reorderBuffer_1_bits_destinationRegister ? io_reorderBuffer_1_bits_value : _GEN_42; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_75 = 5'hb == io_reorderBuffer_1_bits_destinationRegister ? io_reorderBuffer_1_bits_value : _GEN_43; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_76 = 5'hc == io_reorderBuffer_1_bits_destinationRegister ? io_reorderBuffer_1_bits_value : _GEN_44; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_77 = 5'hd == io_reorderBuffer_1_bits_destinationRegister ? io_reorderBuffer_1_bits_value : _GEN_45; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_78 = 5'he == io_reorderBuffer_1_bits_destinationRegister ? io_reorderBuffer_1_bits_value : _GEN_46; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_79 = 5'hf == io_reorderBuffer_1_bits_destinationRegister ? io_reorderBuffer_1_bits_value : _GEN_47; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_80 = 5'h10 == io_reorderBuffer_1_bits_destinationRegister ? io_reorderBuffer_1_bits_value : _GEN_48; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_81 = 5'h11 == io_reorderBuffer_1_bits_destinationRegister ? io_reorderBuffer_1_bits_value : _GEN_49; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_82 = 5'h12 == io_reorderBuffer_1_bits_destinationRegister ? io_reorderBuffer_1_bits_value : _GEN_50; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_83 = 5'h13 == io_reorderBuffer_1_bits_destinationRegister ? io_reorderBuffer_1_bits_value : _GEN_51; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_84 = 5'h14 == io_reorderBuffer_1_bits_destinationRegister ? io_reorderBuffer_1_bits_value : _GEN_52; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_85 = 5'h15 == io_reorderBuffer_1_bits_destinationRegister ? io_reorderBuffer_1_bits_value : _GEN_53; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_86 = 5'h16 == io_reorderBuffer_1_bits_destinationRegister ? io_reorderBuffer_1_bits_value : _GEN_54; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_87 = 5'h17 == io_reorderBuffer_1_bits_destinationRegister ? io_reorderBuffer_1_bits_value : _GEN_55; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_88 = 5'h18 == io_reorderBuffer_1_bits_destinationRegister ? io_reorderBuffer_1_bits_value : _GEN_56; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_89 = 5'h19 == io_reorderBuffer_1_bits_destinationRegister ? io_reorderBuffer_1_bits_value : _GEN_57; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_90 = 5'h1a == io_reorderBuffer_1_bits_destinationRegister ? io_reorderBuffer_1_bits_value : _GEN_58; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_91 = 5'h1b == io_reorderBuffer_1_bits_destinationRegister ? io_reorderBuffer_1_bits_value : _GEN_59; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_92 = 5'h1c == io_reorderBuffer_1_bits_destinationRegister ? io_reorderBuffer_1_bits_value : _GEN_60; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_93 = 5'h1d == io_reorderBuffer_1_bits_destinationRegister ? io_reorderBuffer_1_bits_value : _GEN_61; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_94 = 5'h1e == io_reorderBuffer_1_bits_destinationRegister ? io_reorderBuffer_1_bits_value : _GEN_62; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_95 = 5'h1f == io_reorderBuffer_1_bits_destinationRegister ? io_reorderBuffer_1_bits_value : _GEN_63; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_97 = io_reorderBuffer_1_valid ? _GEN_65 : _GEN_33; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_98 = io_reorderBuffer_1_valid ? _GEN_66 : _GEN_34; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_99 = io_reorderBuffer_1_valid ? _GEN_67 : _GEN_35; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_100 = io_reorderBuffer_1_valid ? _GEN_68 : _GEN_36; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_101 = io_reorderBuffer_1_valid ? _GEN_69 : _GEN_37; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_102 = io_reorderBuffer_1_valid ? _GEN_70 : _GEN_38; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_103 = io_reorderBuffer_1_valid ? _GEN_71 : _GEN_39; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_104 = io_reorderBuffer_1_valid ? _GEN_72 : _GEN_40; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_105 = io_reorderBuffer_1_valid ? _GEN_73 : _GEN_41; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_106 = io_reorderBuffer_1_valid ? _GEN_74 : _GEN_42; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_107 = io_reorderBuffer_1_valid ? _GEN_75 : _GEN_43; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_108 = io_reorderBuffer_1_valid ? _GEN_76 : _GEN_44; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_109 = io_reorderBuffer_1_valid ? _GEN_77 : _GEN_45; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_110 = io_reorderBuffer_1_valid ? _GEN_78 : _GEN_46; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_111 = io_reorderBuffer_1_valid ? _GEN_79 : _GEN_47; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_112 = io_reorderBuffer_1_valid ? _GEN_80 : _GEN_48; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_113 = io_reorderBuffer_1_valid ? _GEN_81 : _GEN_49; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_114 = io_reorderBuffer_1_valid ? _GEN_82 : _GEN_50; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_115 = io_reorderBuffer_1_valid ? _GEN_83 : _GEN_51; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_116 = io_reorderBuffer_1_valid ? _GEN_84 : _GEN_52; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_117 = io_reorderBuffer_1_valid ? _GEN_85 : _GEN_53; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_118 = io_reorderBuffer_1_valid ? _GEN_86 : _GEN_54; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_119 = io_reorderBuffer_1_valid ? _GEN_87 : _GEN_55; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_120 = io_reorderBuffer_1_valid ? _GEN_88 : _GEN_56; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_121 = io_reorderBuffer_1_valid ? _GEN_89 : _GEN_57; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_122 = io_reorderBuffer_1_valid ? _GEN_90 : _GEN_58; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_123 = io_reorderBuffer_1_valid ? _GEN_91 : _GEN_59; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_124 = io_reorderBuffer_1_valid ? _GEN_92 : _GEN_60; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_125 = io_reorderBuffer_1_valid ? _GEN_93 : _GEN_61; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_126 = io_reorderBuffer_1_valid ? _GEN_94 : _GEN_62; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_127 = io_reorderBuffer_1_valid ? _GEN_95 : _GEN_63; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_129 = 5'h1 == io_reorderBuffer_2_bits_destinationRegister ? io_reorderBuffer_2_bits_value : _GEN_97; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_130 = 5'h2 == io_reorderBuffer_2_bits_destinationRegister ? io_reorderBuffer_2_bits_value : _GEN_98; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_131 = 5'h3 == io_reorderBuffer_2_bits_destinationRegister ? io_reorderBuffer_2_bits_value : _GEN_99; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_132 = 5'h4 == io_reorderBuffer_2_bits_destinationRegister ? io_reorderBuffer_2_bits_value : _GEN_100; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_133 = 5'h5 == io_reorderBuffer_2_bits_destinationRegister ? io_reorderBuffer_2_bits_value : _GEN_101; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_134 = 5'h6 == io_reorderBuffer_2_bits_destinationRegister ? io_reorderBuffer_2_bits_value : _GEN_102; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_135 = 5'h7 == io_reorderBuffer_2_bits_destinationRegister ? io_reorderBuffer_2_bits_value : _GEN_103; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_136 = 5'h8 == io_reorderBuffer_2_bits_destinationRegister ? io_reorderBuffer_2_bits_value : _GEN_104; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_137 = 5'h9 == io_reorderBuffer_2_bits_destinationRegister ? io_reorderBuffer_2_bits_value : _GEN_105; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_138 = 5'ha == io_reorderBuffer_2_bits_destinationRegister ? io_reorderBuffer_2_bits_value : _GEN_106; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_139 = 5'hb == io_reorderBuffer_2_bits_destinationRegister ? io_reorderBuffer_2_bits_value : _GEN_107; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_140 = 5'hc == io_reorderBuffer_2_bits_destinationRegister ? io_reorderBuffer_2_bits_value : _GEN_108; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_141 = 5'hd == io_reorderBuffer_2_bits_destinationRegister ? io_reorderBuffer_2_bits_value : _GEN_109; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_142 = 5'he == io_reorderBuffer_2_bits_destinationRegister ? io_reorderBuffer_2_bits_value : _GEN_110; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_143 = 5'hf == io_reorderBuffer_2_bits_destinationRegister ? io_reorderBuffer_2_bits_value : _GEN_111; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_144 = 5'h10 == io_reorderBuffer_2_bits_destinationRegister ? io_reorderBuffer_2_bits_value : _GEN_112
    ; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_145 = 5'h11 == io_reorderBuffer_2_bits_destinationRegister ? io_reorderBuffer_2_bits_value : _GEN_113
    ; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_146 = 5'h12 == io_reorderBuffer_2_bits_destinationRegister ? io_reorderBuffer_2_bits_value : _GEN_114
    ; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_147 = 5'h13 == io_reorderBuffer_2_bits_destinationRegister ? io_reorderBuffer_2_bits_value : _GEN_115
    ; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_148 = 5'h14 == io_reorderBuffer_2_bits_destinationRegister ? io_reorderBuffer_2_bits_value : _GEN_116
    ; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_149 = 5'h15 == io_reorderBuffer_2_bits_destinationRegister ? io_reorderBuffer_2_bits_value : _GEN_117
    ; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_150 = 5'h16 == io_reorderBuffer_2_bits_destinationRegister ? io_reorderBuffer_2_bits_value : _GEN_118
    ; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_151 = 5'h17 == io_reorderBuffer_2_bits_destinationRegister ? io_reorderBuffer_2_bits_value : _GEN_119
    ; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_152 = 5'h18 == io_reorderBuffer_2_bits_destinationRegister ? io_reorderBuffer_2_bits_value : _GEN_120
    ; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_153 = 5'h19 == io_reorderBuffer_2_bits_destinationRegister ? io_reorderBuffer_2_bits_value : _GEN_121
    ; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_154 = 5'h1a == io_reorderBuffer_2_bits_destinationRegister ? io_reorderBuffer_2_bits_value : _GEN_122
    ; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_155 = 5'h1b == io_reorderBuffer_2_bits_destinationRegister ? io_reorderBuffer_2_bits_value : _GEN_123
    ; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_156 = 5'h1c == io_reorderBuffer_2_bits_destinationRegister ? io_reorderBuffer_2_bits_value : _GEN_124
    ; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_157 = 5'h1d == io_reorderBuffer_2_bits_destinationRegister ? io_reorderBuffer_2_bits_value : _GEN_125
    ; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_158 = 5'h1e == io_reorderBuffer_2_bits_destinationRegister ? io_reorderBuffer_2_bits_value : _GEN_126
    ; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_159 = 5'h1f == io_reorderBuffer_2_bits_destinationRegister ? io_reorderBuffer_2_bits_value : _GEN_127
    ; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_161 = io_reorderBuffer_2_valid ? _GEN_129 : _GEN_97; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_162 = io_reorderBuffer_2_valid ? _GEN_130 : _GEN_98; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_163 = io_reorderBuffer_2_valid ? _GEN_131 : _GEN_99; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_164 = io_reorderBuffer_2_valid ? _GEN_132 : _GEN_100; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_165 = io_reorderBuffer_2_valid ? _GEN_133 : _GEN_101; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_166 = io_reorderBuffer_2_valid ? _GEN_134 : _GEN_102; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_167 = io_reorderBuffer_2_valid ? _GEN_135 : _GEN_103; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_168 = io_reorderBuffer_2_valid ? _GEN_136 : _GEN_104; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_169 = io_reorderBuffer_2_valid ? _GEN_137 : _GEN_105; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_170 = io_reorderBuffer_2_valid ? _GEN_138 : _GEN_106; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_171 = io_reorderBuffer_2_valid ? _GEN_139 : _GEN_107; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_172 = io_reorderBuffer_2_valid ? _GEN_140 : _GEN_108; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_173 = io_reorderBuffer_2_valid ? _GEN_141 : _GEN_109; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_174 = io_reorderBuffer_2_valid ? _GEN_142 : _GEN_110; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_175 = io_reorderBuffer_2_valid ? _GEN_143 : _GEN_111; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_176 = io_reorderBuffer_2_valid ? _GEN_144 : _GEN_112; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_177 = io_reorderBuffer_2_valid ? _GEN_145 : _GEN_113; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_178 = io_reorderBuffer_2_valid ? _GEN_146 : _GEN_114; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_179 = io_reorderBuffer_2_valid ? _GEN_147 : _GEN_115; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_180 = io_reorderBuffer_2_valid ? _GEN_148 : _GEN_116; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_181 = io_reorderBuffer_2_valid ? _GEN_149 : _GEN_117; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_182 = io_reorderBuffer_2_valid ? _GEN_150 : _GEN_118; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_183 = io_reorderBuffer_2_valid ? _GEN_151 : _GEN_119; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_184 = io_reorderBuffer_2_valid ? _GEN_152 : _GEN_120; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_185 = io_reorderBuffer_2_valid ? _GEN_153 : _GEN_121; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_186 = io_reorderBuffer_2_valid ? _GEN_154 : _GEN_122; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_187 = io_reorderBuffer_2_valid ? _GEN_155 : _GEN_123; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_188 = io_reorderBuffer_2_valid ? _GEN_156 : _GEN_124; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_189 = io_reorderBuffer_2_valid ? _GEN_157 : _GEN_125; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_190 = io_reorderBuffer_2_valid ? _GEN_158 : _GEN_126; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_191 = io_reorderBuffer_2_valid ? _GEN_159 : _GEN_127; // @[RegisterFile.scala 45:20]
  wire  _io_decoders_0_value1_T = io_decoders_0_sourceRegister1 == 5'h0; // @[RegisterFile.scala 54:27]
  wire [63:0] _GEN_257 = 5'h1 == io_decoders_0_sourceRegister1 ? registers_1 : 64'h0; // @[RegisterFile.scala 53:{22,22}]
  wire [63:0] _GEN_258 = 5'h2 == io_decoders_0_sourceRegister1 ? registers_2 : _GEN_257; // @[RegisterFile.scala 53:{22,22}]
  wire [63:0] _GEN_259 = 5'h3 == io_decoders_0_sourceRegister1 ? registers_3 : _GEN_258; // @[RegisterFile.scala 53:{22,22}]
  wire [63:0] _GEN_260 = 5'h4 == io_decoders_0_sourceRegister1 ? registers_4 : _GEN_259; // @[RegisterFile.scala 53:{22,22}]
  wire [63:0] _GEN_261 = 5'h5 == io_decoders_0_sourceRegister1 ? registers_5 : _GEN_260; // @[RegisterFile.scala 53:{22,22}]
  wire [63:0] _GEN_262 = 5'h6 == io_decoders_0_sourceRegister1 ? registers_6 : _GEN_261; // @[RegisterFile.scala 53:{22,22}]
  wire [63:0] _GEN_263 = 5'h7 == io_decoders_0_sourceRegister1 ? registers_7 : _GEN_262; // @[RegisterFile.scala 53:{22,22}]
  wire [63:0] _GEN_264 = 5'h8 == io_decoders_0_sourceRegister1 ? registers_8 : _GEN_263; // @[RegisterFile.scala 53:{22,22}]
  wire [63:0] _GEN_265 = 5'h9 == io_decoders_0_sourceRegister1 ? registers_9 : _GEN_264; // @[RegisterFile.scala 53:{22,22}]
  wire [63:0] _GEN_266 = 5'ha == io_decoders_0_sourceRegister1 ? registers_10 : _GEN_265; // @[RegisterFile.scala 53:{22,22}]
  wire [63:0] _GEN_267 = 5'hb == io_decoders_0_sourceRegister1 ? registers_11 : _GEN_266; // @[RegisterFile.scala 53:{22,22}]
  wire [63:0] _GEN_268 = 5'hc == io_decoders_0_sourceRegister1 ? registers_12 : _GEN_267; // @[RegisterFile.scala 53:{22,22}]
  wire [63:0] _GEN_269 = 5'hd == io_decoders_0_sourceRegister1 ? registers_13 : _GEN_268; // @[RegisterFile.scala 53:{22,22}]
  wire [63:0] _GEN_270 = 5'he == io_decoders_0_sourceRegister1 ? registers_14 : _GEN_269; // @[RegisterFile.scala 53:{22,22}]
  wire [63:0] _GEN_271 = 5'hf == io_decoders_0_sourceRegister1 ? registers_15 : _GEN_270; // @[RegisterFile.scala 53:{22,22}]
  wire [63:0] _GEN_272 = 5'h10 == io_decoders_0_sourceRegister1 ? registers_16 : _GEN_271; // @[RegisterFile.scala 53:{22,22}]
  wire [63:0] _GEN_273 = 5'h11 == io_decoders_0_sourceRegister1 ? registers_17 : _GEN_272; // @[RegisterFile.scala 53:{22,22}]
  wire [63:0] _GEN_274 = 5'h12 == io_decoders_0_sourceRegister1 ? registers_18 : _GEN_273; // @[RegisterFile.scala 53:{22,22}]
  wire [63:0] _GEN_275 = 5'h13 == io_decoders_0_sourceRegister1 ? registers_19 : _GEN_274; // @[RegisterFile.scala 53:{22,22}]
  wire [63:0] _GEN_276 = 5'h14 == io_decoders_0_sourceRegister1 ? registers_20 : _GEN_275; // @[RegisterFile.scala 53:{22,22}]
  wire [63:0] _GEN_277 = 5'h15 == io_decoders_0_sourceRegister1 ? registers_21 : _GEN_276; // @[RegisterFile.scala 53:{22,22}]
  wire [63:0] _GEN_278 = 5'h16 == io_decoders_0_sourceRegister1 ? registers_22 : _GEN_277; // @[RegisterFile.scala 53:{22,22}]
  wire [63:0] _GEN_279 = 5'h17 == io_decoders_0_sourceRegister1 ? registers_23 : _GEN_278; // @[RegisterFile.scala 53:{22,22}]
  wire [63:0] _GEN_280 = 5'h18 == io_decoders_0_sourceRegister1 ? registers_24 : _GEN_279; // @[RegisterFile.scala 53:{22,22}]
  wire [63:0] _GEN_281 = 5'h19 == io_decoders_0_sourceRegister1 ? registers_25 : _GEN_280; // @[RegisterFile.scala 53:{22,22}]
  wire [63:0] _GEN_282 = 5'h1a == io_decoders_0_sourceRegister1 ? registers_26 : _GEN_281; // @[RegisterFile.scala 53:{22,22}]
  wire [63:0] _GEN_283 = 5'h1b == io_decoders_0_sourceRegister1 ? registers_27 : _GEN_282; // @[RegisterFile.scala 53:{22,22}]
  wire [63:0] _GEN_284 = 5'h1c == io_decoders_0_sourceRegister1 ? registers_28 : _GEN_283; // @[RegisterFile.scala 53:{22,22}]
  wire [63:0] _GEN_285 = 5'h1d == io_decoders_0_sourceRegister1 ? registers_29 : _GEN_284; // @[RegisterFile.scala 53:{22,22}]
  wire [63:0] _GEN_286 = 5'h1e == io_decoders_0_sourceRegister1 ? registers_30 : _GEN_285; // @[RegisterFile.scala 53:{22,22}]
  wire [63:0] _GEN_287 = 5'h1f == io_decoders_0_sourceRegister1 ? registers_31 : _GEN_286; // @[RegisterFile.scala 53:{22,22}]
  wire  _io_decoders_0_value2_T = io_decoders_0_sourceRegister2 == 5'h0; // @[RegisterFile.scala 59:27]
  wire [63:0] _GEN_289 = 5'h1 == io_decoders_0_sourceRegister2 ? registers_1 : 64'h0; // @[RegisterFile.scala 58:{22,22}]
  wire [63:0] _GEN_290 = 5'h2 == io_decoders_0_sourceRegister2 ? registers_2 : _GEN_289; // @[RegisterFile.scala 58:{22,22}]
  wire [63:0] _GEN_291 = 5'h3 == io_decoders_0_sourceRegister2 ? registers_3 : _GEN_290; // @[RegisterFile.scala 58:{22,22}]
  wire [63:0] _GEN_292 = 5'h4 == io_decoders_0_sourceRegister2 ? registers_4 : _GEN_291; // @[RegisterFile.scala 58:{22,22}]
  wire [63:0] _GEN_293 = 5'h5 == io_decoders_0_sourceRegister2 ? registers_5 : _GEN_292; // @[RegisterFile.scala 58:{22,22}]
  wire [63:0] _GEN_294 = 5'h6 == io_decoders_0_sourceRegister2 ? registers_6 : _GEN_293; // @[RegisterFile.scala 58:{22,22}]
  wire [63:0] _GEN_295 = 5'h7 == io_decoders_0_sourceRegister2 ? registers_7 : _GEN_294; // @[RegisterFile.scala 58:{22,22}]
  wire [63:0] _GEN_296 = 5'h8 == io_decoders_0_sourceRegister2 ? registers_8 : _GEN_295; // @[RegisterFile.scala 58:{22,22}]
  wire [63:0] _GEN_297 = 5'h9 == io_decoders_0_sourceRegister2 ? registers_9 : _GEN_296; // @[RegisterFile.scala 58:{22,22}]
  wire [63:0] _GEN_298 = 5'ha == io_decoders_0_sourceRegister2 ? registers_10 : _GEN_297; // @[RegisterFile.scala 58:{22,22}]
  wire [63:0] _GEN_299 = 5'hb == io_decoders_0_sourceRegister2 ? registers_11 : _GEN_298; // @[RegisterFile.scala 58:{22,22}]
  wire [63:0] _GEN_300 = 5'hc == io_decoders_0_sourceRegister2 ? registers_12 : _GEN_299; // @[RegisterFile.scala 58:{22,22}]
  wire [63:0] _GEN_301 = 5'hd == io_decoders_0_sourceRegister2 ? registers_13 : _GEN_300; // @[RegisterFile.scala 58:{22,22}]
  wire [63:0] _GEN_302 = 5'he == io_decoders_0_sourceRegister2 ? registers_14 : _GEN_301; // @[RegisterFile.scala 58:{22,22}]
  wire [63:0] _GEN_303 = 5'hf == io_decoders_0_sourceRegister2 ? registers_15 : _GEN_302; // @[RegisterFile.scala 58:{22,22}]
  wire [63:0] _GEN_304 = 5'h10 == io_decoders_0_sourceRegister2 ? registers_16 : _GEN_303; // @[RegisterFile.scala 58:{22,22}]
  wire [63:0] _GEN_305 = 5'h11 == io_decoders_0_sourceRegister2 ? registers_17 : _GEN_304; // @[RegisterFile.scala 58:{22,22}]
  wire [63:0] _GEN_306 = 5'h12 == io_decoders_0_sourceRegister2 ? registers_18 : _GEN_305; // @[RegisterFile.scala 58:{22,22}]
  wire [63:0] _GEN_307 = 5'h13 == io_decoders_0_sourceRegister2 ? registers_19 : _GEN_306; // @[RegisterFile.scala 58:{22,22}]
  wire [63:0] _GEN_308 = 5'h14 == io_decoders_0_sourceRegister2 ? registers_20 : _GEN_307; // @[RegisterFile.scala 58:{22,22}]
  wire [63:0] _GEN_309 = 5'h15 == io_decoders_0_sourceRegister2 ? registers_21 : _GEN_308; // @[RegisterFile.scala 58:{22,22}]
  wire [63:0] _GEN_310 = 5'h16 == io_decoders_0_sourceRegister2 ? registers_22 : _GEN_309; // @[RegisterFile.scala 58:{22,22}]
  wire [63:0] _GEN_311 = 5'h17 == io_decoders_0_sourceRegister2 ? registers_23 : _GEN_310; // @[RegisterFile.scala 58:{22,22}]
  wire [63:0] _GEN_312 = 5'h18 == io_decoders_0_sourceRegister2 ? registers_24 : _GEN_311; // @[RegisterFile.scala 58:{22,22}]
  wire [63:0] _GEN_313 = 5'h19 == io_decoders_0_sourceRegister2 ? registers_25 : _GEN_312; // @[RegisterFile.scala 58:{22,22}]
  wire [63:0] _GEN_314 = 5'h1a == io_decoders_0_sourceRegister2 ? registers_26 : _GEN_313; // @[RegisterFile.scala 58:{22,22}]
  wire [63:0] _GEN_315 = 5'h1b == io_decoders_0_sourceRegister2 ? registers_27 : _GEN_314; // @[RegisterFile.scala 58:{22,22}]
  wire [63:0] _GEN_316 = 5'h1c == io_decoders_0_sourceRegister2 ? registers_28 : _GEN_315; // @[RegisterFile.scala 58:{22,22}]
  wire [63:0] _GEN_317 = 5'h1d == io_decoders_0_sourceRegister2 ? registers_29 : _GEN_316; // @[RegisterFile.scala 58:{22,22}]
  wire [63:0] _GEN_318 = 5'h1e == io_decoders_0_sourceRegister2 ? registers_30 : _GEN_317; // @[RegisterFile.scala 58:{22,22}]
  wire [63:0] _GEN_319 = 5'h1f == io_decoders_0_sourceRegister2 ? registers_31 : _GEN_318; // @[RegisterFile.scala 58:{22,22}]
  assign io_decoders_0_value1 = _io_decoders_0_value1_T ? 64'h0 : _GEN_287; // @[RegisterFile.scala 53:22]
  assign io_decoders_0_value2 = _io_decoders_0_value2_T ? 64'h0 : _GEN_319; // @[RegisterFile.scala 58:22]
  always @(posedge clock) begin
    if (reset) begin // @[RegisterFile.scala 37:26]
      registers_1 <= 64'h0; // @[RegisterFile.scala 37:26]
    end else if (io_reorderBuffer_3_valid) begin // @[RegisterFile.scala 45:20]
      if (5'h1 == io_reorderBuffer_3_bits_destinationRegister) begin // @[RegisterFile.scala 46:46]
        registers_1 <= io_reorderBuffer_3_bits_value; // @[RegisterFile.scala 46:46]
      end else begin
        registers_1 <= _GEN_161;
      end
    end else begin
      registers_1 <= _GEN_161;
    end
    if (reset) begin // @[RegisterFile.scala 37:26]
      registers_2 <= 64'h0; // @[RegisterFile.scala 37:26]
    end else if (io_reorderBuffer_3_valid) begin // @[RegisterFile.scala 45:20]
      if (5'h2 == io_reorderBuffer_3_bits_destinationRegister) begin // @[RegisterFile.scala 46:46]
        registers_2 <= io_reorderBuffer_3_bits_value; // @[RegisterFile.scala 46:46]
      end else begin
        registers_2 <= _GEN_162;
      end
    end else begin
      registers_2 <= _GEN_162;
    end
    if (reset) begin // @[RegisterFile.scala 37:26]
      registers_3 <= 64'h0; // @[RegisterFile.scala 37:26]
    end else if (io_reorderBuffer_3_valid) begin // @[RegisterFile.scala 45:20]
      if (5'h3 == io_reorderBuffer_3_bits_destinationRegister) begin // @[RegisterFile.scala 46:46]
        registers_3 <= io_reorderBuffer_3_bits_value; // @[RegisterFile.scala 46:46]
      end else begin
        registers_3 <= _GEN_163;
      end
    end else begin
      registers_3 <= _GEN_163;
    end
    if (reset) begin // @[RegisterFile.scala 37:26]
      registers_4 <= 64'h0; // @[RegisterFile.scala 37:26]
    end else if (io_reorderBuffer_3_valid) begin // @[RegisterFile.scala 45:20]
      if (5'h4 == io_reorderBuffer_3_bits_destinationRegister) begin // @[RegisterFile.scala 46:46]
        registers_4 <= io_reorderBuffer_3_bits_value; // @[RegisterFile.scala 46:46]
      end else begin
        registers_4 <= _GEN_164;
      end
    end else begin
      registers_4 <= _GEN_164;
    end
    if (reset) begin // @[RegisterFile.scala 37:26]
      registers_5 <= 64'h0; // @[RegisterFile.scala 37:26]
    end else if (io_reorderBuffer_3_valid) begin // @[RegisterFile.scala 45:20]
      if (5'h5 == io_reorderBuffer_3_bits_destinationRegister) begin // @[RegisterFile.scala 46:46]
        registers_5 <= io_reorderBuffer_3_bits_value; // @[RegisterFile.scala 46:46]
      end else begin
        registers_5 <= _GEN_165;
      end
    end else begin
      registers_5 <= _GEN_165;
    end
    if (reset) begin // @[RegisterFile.scala 37:26]
      registers_6 <= 64'h0; // @[RegisterFile.scala 37:26]
    end else if (io_reorderBuffer_3_valid) begin // @[RegisterFile.scala 45:20]
      if (5'h6 == io_reorderBuffer_3_bits_destinationRegister) begin // @[RegisterFile.scala 46:46]
        registers_6 <= io_reorderBuffer_3_bits_value; // @[RegisterFile.scala 46:46]
      end else begin
        registers_6 <= _GEN_166;
      end
    end else begin
      registers_6 <= _GEN_166;
    end
    if (reset) begin // @[RegisterFile.scala 37:26]
      registers_7 <= 64'h0; // @[RegisterFile.scala 37:26]
    end else if (io_reorderBuffer_3_valid) begin // @[RegisterFile.scala 45:20]
      if (5'h7 == io_reorderBuffer_3_bits_destinationRegister) begin // @[RegisterFile.scala 46:46]
        registers_7 <= io_reorderBuffer_3_bits_value; // @[RegisterFile.scala 46:46]
      end else begin
        registers_7 <= _GEN_167;
      end
    end else begin
      registers_7 <= _GEN_167;
    end
    if (reset) begin // @[RegisterFile.scala 37:26]
      registers_8 <= 64'h0; // @[RegisterFile.scala 37:26]
    end else if (io_reorderBuffer_3_valid) begin // @[RegisterFile.scala 45:20]
      if (5'h8 == io_reorderBuffer_3_bits_destinationRegister) begin // @[RegisterFile.scala 46:46]
        registers_8 <= io_reorderBuffer_3_bits_value; // @[RegisterFile.scala 46:46]
      end else begin
        registers_8 <= _GEN_168;
      end
    end else begin
      registers_8 <= _GEN_168;
    end
    if (reset) begin // @[RegisterFile.scala 37:26]
      registers_9 <= 64'h0; // @[RegisterFile.scala 37:26]
    end else if (io_reorderBuffer_3_valid) begin // @[RegisterFile.scala 45:20]
      if (5'h9 == io_reorderBuffer_3_bits_destinationRegister) begin // @[RegisterFile.scala 46:46]
        registers_9 <= io_reorderBuffer_3_bits_value; // @[RegisterFile.scala 46:46]
      end else begin
        registers_9 <= _GEN_169;
      end
    end else begin
      registers_9 <= _GEN_169;
    end
    if (reset) begin // @[RegisterFile.scala 37:26]
      registers_10 <= 64'h0; // @[RegisterFile.scala 37:26]
    end else if (io_reorderBuffer_3_valid) begin // @[RegisterFile.scala 45:20]
      if (5'ha == io_reorderBuffer_3_bits_destinationRegister) begin // @[RegisterFile.scala 46:46]
        registers_10 <= io_reorderBuffer_3_bits_value; // @[RegisterFile.scala 46:46]
      end else begin
        registers_10 <= _GEN_170;
      end
    end else begin
      registers_10 <= _GEN_170;
    end
    if (reset) begin // @[RegisterFile.scala 37:26]
      registers_11 <= 64'h0; // @[RegisterFile.scala 37:26]
    end else if (io_reorderBuffer_3_valid) begin // @[RegisterFile.scala 45:20]
      if (5'hb == io_reorderBuffer_3_bits_destinationRegister) begin // @[RegisterFile.scala 46:46]
        registers_11 <= io_reorderBuffer_3_bits_value; // @[RegisterFile.scala 46:46]
      end else begin
        registers_11 <= _GEN_171;
      end
    end else begin
      registers_11 <= _GEN_171;
    end
    if (reset) begin // @[RegisterFile.scala 37:26]
      registers_12 <= 64'h0; // @[RegisterFile.scala 37:26]
    end else if (io_reorderBuffer_3_valid) begin // @[RegisterFile.scala 45:20]
      if (5'hc == io_reorderBuffer_3_bits_destinationRegister) begin // @[RegisterFile.scala 46:46]
        registers_12 <= io_reorderBuffer_3_bits_value; // @[RegisterFile.scala 46:46]
      end else begin
        registers_12 <= _GEN_172;
      end
    end else begin
      registers_12 <= _GEN_172;
    end
    if (reset) begin // @[RegisterFile.scala 37:26]
      registers_13 <= 64'h0; // @[RegisterFile.scala 37:26]
    end else if (io_reorderBuffer_3_valid) begin // @[RegisterFile.scala 45:20]
      if (5'hd == io_reorderBuffer_3_bits_destinationRegister) begin // @[RegisterFile.scala 46:46]
        registers_13 <= io_reorderBuffer_3_bits_value; // @[RegisterFile.scala 46:46]
      end else begin
        registers_13 <= _GEN_173;
      end
    end else begin
      registers_13 <= _GEN_173;
    end
    if (reset) begin // @[RegisterFile.scala 37:26]
      registers_14 <= 64'h0; // @[RegisterFile.scala 37:26]
    end else if (io_reorderBuffer_3_valid) begin // @[RegisterFile.scala 45:20]
      if (5'he == io_reorderBuffer_3_bits_destinationRegister) begin // @[RegisterFile.scala 46:46]
        registers_14 <= io_reorderBuffer_3_bits_value; // @[RegisterFile.scala 46:46]
      end else begin
        registers_14 <= _GEN_174;
      end
    end else begin
      registers_14 <= _GEN_174;
    end
    if (reset) begin // @[RegisterFile.scala 37:26]
      registers_15 <= 64'h0; // @[RegisterFile.scala 37:26]
    end else if (io_reorderBuffer_3_valid) begin // @[RegisterFile.scala 45:20]
      if (5'hf == io_reorderBuffer_3_bits_destinationRegister) begin // @[RegisterFile.scala 46:46]
        registers_15 <= io_reorderBuffer_3_bits_value; // @[RegisterFile.scala 46:46]
      end else begin
        registers_15 <= _GEN_175;
      end
    end else begin
      registers_15 <= _GEN_175;
    end
    if (reset) begin // @[RegisterFile.scala 37:26]
      registers_16 <= 64'h0; // @[RegisterFile.scala 37:26]
    end else if (io_reorderBuffer_3_valid) begin // @[RegisterFile.scala 45:20]
      if (5'h10 == io_reorderBuffer_3_bits_destinationRegister) begin // @[RegisterFile.scala 46:46]
        registers_16 <= io_reorderBuffer_3_bits_value; // @[RegisterFile.scala 46:46]
      end else begin
        registers_16 <= _GEN_176;
      end
    end else begin
      registers_16 <= _GEN_176;
    end
    if (reset) begin // @[RegisterFile.scala 37:26]
      registers_17 <= 64'h0; // @[RegisterFile.scala 37:26]
    end else if (io_reorderBuffer_3_valid) begin // @[RegisterFile.scala 45:20]
      if (5'h11 == io_reorderBuffer_3_bits_destinationRegister) begin // @[RegisterFile.scala 46:46]
        registers_17 <= io_reorderBuffer_3_bits_value; // @[RegisterFile.scala 46:46]
      end else begin
        registers_17 <= _GEN_177;
      end
    end else begin
      registers_17 <= _GEN_177;
    end
    if (reset) begin // @[RegisterFile.scala 37:26]
      registers_18 <= 64'h0; // @[RegisterFile.scala 37:26]
    end else if (io_reorderBuffer_3_valid) begin // @[RegisterFile.scala 45:20]
      if (5'h12 == io_reorderBuffer_3_bits_destinationRegister) begin // @[RegisterFile.scala 46:46]
        registers_18 <= io_reorderBuffer_3_bits_value; // @[RegisterFile.scala 46:46]
      end else begin
        registers_18 <= _GEN_178;
      end
    end else begin
      registers_18 <= _GEN_178;
    end
    if (reset) begin // @[RegisterFile.scala 37:26]
      registers_19 <= 64'h0; // @[RegisterFile.scala 37:26]
    end else if (io_reorderBuffer_3_valid) begin // @[RegisterFile.scala 45:20]
      if (5'h13 == io_reorderBuffer_3_bits_destinationRegister) begin // @[RegisterFile.scala 46:46]
        registers_19 <= io_reorderBuffer_3_bits_value; // @[RegisterFile.scala 46:46]
      end else begin
        registers_19 <= _GEN_179;
      end
    end else begin
      registers_19 <= _GEN_179;
    end
    if (reset) begin // @[RegisterFile.scala 37:26]
      registers_20 <= 64'h0; // @[RegisterFile.scala 37:26]
    end else if (io_reorderBuffer_3_valid) begin // @[RegisterFile.scala 45:20]
      if (5'h14 == io_reorderBuffer_3_bits_destinationRegister) begin // @[RegisterFile.scala 46:46]
        registers_20 <= io_reorderBuffer_3_bits_value; // @[RegisterFile.scala 46:46]
      end else begin
        registers_20 <= _GEN_180;
      end
    end else begin
      registers_20 <= _GEN_180;
    end
    if (reset) begin // @[RegisterFile.scala 37:26]
      registers_21 <= 64'h0; // @[RegisterFile.scala 37:26]
    end else if (io_reorderBuffer_3_valid) begin // @[RegisterFile.scala 45:20]
      if (5'h15 == io_reorderBuffer_3_bits_destinationRegister) begin // @[RegisterFile.scala 46:46]
        registers_21 <= io_reorderBuffer_3_bits_value; // @[RegisterFile.scala 46:46]
      end else begin
        registers_21 <= _GEN_181;
      end
    end else begin
      registers_21 <= _GEN_181;
    end
    if (reset) begin // @[RegisterFile.scala 37:26]
      registers_22 <= 64'h0; // @[RegisterFile.scala 37:26]
    end else if (io_reorderBuffer_3_valid) begin // @[RegisterFile.scala 45:20]
      if (5'h16 == io_reorderBuffer_3_bits_destinationRegister) begin // @[RegisterFile.scala 46:46]
        registers_22 <= io_reorderBuffer_3_bits_value; // @[RegisterFile.scala 46:46]
      end else begin
        registers_22 <= _GEN_182;
      end
    end else begin
      registers_22 <= _GEN_182;
    end
    if (reset) begin // @[RegisterFile.scala 37:26]
      registers_23 <= 64'h0; // @[RegisterFile.scala 37:26]
    end else if (io_reorderBuffer_3_valid) begin // @[RegisterFile.scala 45:20]
      if (5'h17 == io_reorderBuffer_3_bits_destinationRegister) begin // @[RegisterFile.scala 46:46]
        registers_23 <= io_reorderBuffer_3_bits_value; // @[RegisterFile.scala 46:46]
      end else begin
        registers_23 <= _GEN_183;
      end
    end else begin
      registers_23 <= _GEN_183;
    end
    if (reset) begin // @[RegisterFile.scala 37:26]
      registers_24 <= 64'h0; // @[RegisterFile.scala 37:26]
    end else if (io_reorderBuffer_3_valid) begin // @[RegisterFile.scala 45:20]
      if (5'h18 == io_reorderBuffer_3_bits_destinationRegister) begin // @[RegisterFile.scala 46:46]
        registers_24 <= io_reorderBuffer_3_bits_value; // @[RegisterFile.scala 46:46]
      end else begin
        registers_24 <= _GEN_184;
      end
    end else begin
      registers_24 <= _GEN_184;
    end
    if (reset) begin // @[RegisterFile.scala 37:26]
      registers_25 <= 64'h0; // @[RegisterFile.scala 37:26]
    end else if (io_reorderBuffer_3_valid) begin // @[RegisterFile.scala 45:20]
      if (5'h19 == io_reorderBuffer_3_bits_destinationRegister) begin // @[RegisterFile.scala 46:46]
        registers_25 <= io_reorderBuffer_3_bits_value; // @[RegisterFile.scala 46:46]
      end else begin
        registers_25 <= _GEN_185;
      end
    end else begin
      registers_25 <= _GEN_185;
    end
    if (reset) begin // @[RegisterFile.scala 37:26]
      registers_26 <= 64'h0; // @[RegisterFile.scala 37:26]
    end else if (io_reorderBuffer_3_valid) begin // @[RegisterFile.scala 45:20]
      if (5'h1a == io_reorderBuffer_3_bits_destinationRegister) begin // @[RegisterFile.scala 46:46]
        registers_26 <= io_reorderBuffer_3_bits_value; // @[RegisterFile.scala 46:46]
      end else begin
        registers_26 <= _GEN_186;
      end
    end else begin
      registers_26 <= _GEN_186;
    end
    if (reset) begin // @[RegisterFile.scala 37:26]
      registers_27 <= 64'h0; // @[RegisterFile.scala 37:26]
    end else if (io_reorderBuffer_3_valid) begin // @[RegisterFile.scala 45:20]
      if (5'h1b == io_reorderBuffer_3_bits_destinationRegister) begin // @[RegisterFile.scala 46:46]
        registers_27 <= io_reorderBuffer_3_bits_value; // @[RegisterFile.scala 46:46]
      end else begin
        registers_27 <= _GEN_187;
      end
    end else begin
      registers_27 <= _GEN_187;
    end
    if (reset) begin // @[RegisterFile.scala 37:26]
      registers_28 <= 64'h0; // @[RegisterFile.scala 37:26]
    end else if (io_reorderBuffer_3_valid) begin // @[RegisterFile.scala 45:20]
      if (5'h1c == io_reorderBuffer_3_bits_destinationRegister) begin // @[RegisterFile.scala 46:46]
        registers_28 <= io_reorderBuffer_3_bits_value; // @[RegisterFile.scala 46:46]
      end else begin
        registers_28 <= _GEN_188;
      end
    end else begin
      registers_28 <= _GEN_188;
    end
    if (reset) begin // @[RegisterFile.scala 37:26]
      registers_29 <= 64'h0; // @[RegisterFile.scala 37:26]
    end else if (io_reorderBuffer_3_valid) begin // @[RegisterFile.scala 45:20]
      if (5'h1d == io_reorderBuffer_3_bits_destinationRegister) begin // @[RegisterFile.scala 46:46]
        registers_29 <= io_reorderBuffer_3_bits_value; // @[RegisterFile.scala 46:46]
      end else begin
        registers_29 <= _GEN_189;
      end
    end else begin
      registers_29 <= _GEN_189;
    end
    if (reset) begin // @[RegisterFile.scala 37:26]
      registers_30 <= 64'h0; // @[RegisterFile.scala 37:26]
    end else if (io_reorderBuffer_3_valid) begin // @[RegisterFile.scala 45:20]
      if (5'h1e == io_reorderBuffer_3_bits_destinationRegister) begin // @[RegisterFile.scala 46:46]
        registers_30 <= io_reorderBuffer_3_bits_value; // @[RegisterFile.scala 46:46]
      end else begin
        registers_30 <= _GEN_190;
      end
    end else begin
      registers_30 <= _GEN_190;
    end
    if (reset) begin // @[RegisterFile.scala 37:26]
      registers_31 <= 64'h0; // @[RegisterFile.scala 37:26]
    end else if (io_reorderBuffer_3_valid) begin // @[RegisterFile.scala 45:20]
      if (5'h1f == io_reorderBuffer_3_bits_destinationRegister) begin // @[RegisterFile.scala 46:46]
        registers_31 <= io_reorderBuffer_3_bits_value; // @[RegisterFile.scala 46:46]
      end else begin
        registers_31 <= _GEN_191;
      end
    end else begin
      registers_31 <= _GEN_191;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  registers_1 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  registers_2 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  registers_3 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  registers_4 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  registers_5 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  registers_6 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  registers_7 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  registers_8 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  registers_9 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  registers_10 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  registers_11 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  registers_12 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  registers_13 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  registers_14 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  registers_15 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  registers_16 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  registers_17 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  registers_18 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  registers_19 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  registers_20 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  registers_21 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  registers_22 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  registers_23 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  registers_24 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  registers_25 = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  registers_26 = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  registers_27 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  registers_28 = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  registers_29 = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  registers_30 = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  registers_31 = _RAND_30[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RegisterFile_1(
  input         clock,
  input         reset,
  input  [4:0]  io_decoders_0_sourceRegister1,
  input  [4:0]  io_decoders_0_sourceRegister2,
  output [63:0] io_decoders_0_value1,
  output [63:0] io_decoders_0_value2,
  input         io_reorderBuffer_0_valid,
  input  [4:0]  io_reorderBuffer_0_bits_destinationRegister,
  input  [63:0] io_reorderBuffer_0_bits_value,
  input         io_reorderBuffer_1_valid,
  input  [4:0]  io_reorderBuffer_1_bits_destinationRegister,
  input  [63:0] io_reorderBuffer_1_bits_value,
  input         io_reorderBuffer_2_valid,
  input  [4:0]  io_reorderBuffer_2_bits_destinationRegister,
  input  [63:0] io_reorderBuffer_2_bits_value,
  input         io_reorderBuffer_3_valid,
  input  [4:0]  io_reorderBuffer_3_bits_destinationRegister,
  input  [63:0] io_reorderBuffer_3_bits_value
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] registers_1; // @[RegisterFile.scala 37:26]
  reg [63:0] registers_2; // @[RegisterFile.scala 37:26]
  reg [63:0] registers_3; // @[RegisterFile.scala 37:26]
  reg [63:0] registers_4; // @[RegisterFile.scala 37:26]
  reg [63:0] registers_5; // @[RegisterFile.scala 37:26]
  reg [63:0] registers_6; // @[RegisterFile.scala 37:26]
  reg [63:0] registers_7; // @[RegisterFile.scala 37:26]
  reg [63:0] registers_8; // @[RegisterFile.scala 37:26]
  reg [63:0] registers_9; // @[RegisterFile.scala 37:26]
  reg [63:0] registers_10; // @[RegisterFile.scala 37:26]
  reg [63:0] registers_11; // @[RegisterFile.scala 37:26]
  reg [63:0] registers_12; // @[RegisterFile.scala 37:26]
  reg [63:0] registers_13; // @[RegisterFile.scala 37:26]
  reg [63:0] registers_14; // @[RegisterFile.scala 37:26]
  reg [63:0] registers_15; // @[RegisterFile.scala 37:26]
  reg [63:0] registers_16; // @[RegisterFile.scala 37:26]
  reg [63:0] registers_17; // @[RegisterFile.scala 37:26]
  reg [63:0] registers_18; // @[RegisterFile.scala 37:26]
  reg [63:0] registers_19; // @[RegisterFile.scala 37:26]
  reg [63:0] registers_20; // @[RegisterFile.scala 37:26]
  reg [63:0] registers_21; // @[RegisterFile.scala 37:26]
  reg [63:0] registers_22; // @[RegisterFile.scala 37:26]
  reg [63:0] registers_23; // @[RegisterFile.scala 37:26]
  reg [63:0] registers_24; // @[RegisterFile.scala 37:26]
  reg [63:0] registers_25; // @[RegisterFile.scala 37:26]
  reg [63:0] registers_26; // @[RegisterFile.scala 37:26]
  reg [63:0] registers_27; // @[RegisterFile.scala 37:26]
  reg [63:0] registers_28; // @[RegisterFile.scala 37:26]
  reg [63:0] registers_29; // @[RegisterFile.scala 37:26]
  reg [63:0] registers_30; // @[RegisterFile.scala 37:26]
  reg [63:0] registers_31; // @[RegisterFile.scala 37:26]
  wire [63:0] _GEN_1 = 5'h1 == io_reorderBuffer_0_bits_destinationRegister ? io_reorderBuffer_0_bits_value : registers_1
    ; // @[RegisterFile.scala 37:26 46:{46,46}]
  wire [63:0] _GEN_2 = 5'h2 == io_reorderBuffer_0_bits_destinationRegister ? io_reorderBuffer_0_bits_value : registers_2
    ; // @[RegisterFile.scala 37:26 46:{46,46}]
  wire [63:0] _GEN_3 = 5'h3 == io_reorderBuffer_0_bits_destinationRegister ? io_reorderBuffer_0_bits_value : registers_3
    ; // @[RegisterFile.scala 37:26 46:{46,46}]
  wire [63:0] _GEN_4 = 5'h4 == io_reorderBuffer_0_bits_destinationRegister ? io_reorderBuffer_0_bits_value : registers_4
    ; // @[RegisterFile.scala 37:26 46:{46,46}]
  wire [63:0] _GEN_5 = 5'h5 == io_reorderBuffer_0_bits_destinationRegister ? io_reorderBuffer_0_bits_value : registers_5
    ; // @[RegisterFile.scala 37:26 46:{46,46}]
  wire [63:0] _GEN_6 = 5'h6 == io_reorderBuffer_0_bits_destinationRegister ? io_reorderBuffer_0_bits_value : registers_6
    ; // @[RegisterFile.scala 37:26 46:{46,46}]
  wire [63:0] _GEN_7 = 5'h7 == io_reorderBuffer_0_bits_destinationRegister ? io_reorderBuffer_0_bits_value : registers_7
    ; // @[RegisterFile.scala 37:26 46:{46,46}]
  wire [63:0] _GEN_8 = 5'h8 == io_reorderBuffer_0_bits_destinationRegister ? io_reorderBuffer_0_bits_value : registers_8
    ; // @[RegisterFile.scala 37:26 46:{46,46}]
  wire [63:0] _GEN_9 = 5'h9 == io_reorderBuffer_0_bits_destinationRegister ? io_reorderBuffer_0_bits_value : registers_9
    ; // @[RegisterFile.scala 37:26 46:{46,46}]
  wire [63:0] _GEN_10 = 5'ha == io_reorderBuffer_0_bits_destinationRegister ? io_reorderBuffer_0_bits_value :
    registers_10; // @[RegisterFile.scala 37:26 46:{46,46}]
  wire [63:0] _GEN_11 = 5'hb == io_reorderBuffer_0_bits_destinationRegister ? io_reorderBuffer_0_bits_value :
    registers_11; // @[RegisterFile.scala 37:26 46:{46,46}]
  wire [63:0] _GEN_12 = 5'hc == io_reorderBuffer_0_bits_destinationRegister ? io_reorderBuffer_0_bits_value :
    registers_12; // @[RegisterFile.scala 37:26 46:{46,46}]
  wire [63:0] _GEN_13 = 5'hd == io_reorderBuffer_0_bits_destinationRegister ? io_reorderBuffer_0_bits_value :
    registers_13; // @[RegisterFile.scala 37:26 46:{46,46}]
  wire [63:0] _GEN_14 = 5'he == io_reorderBuffer_0_bits_destinationRegister ? io_reorderBuffer_0_bits_value :
    registers_14; // @[RegisterFile.scala 37:26 46:{46,46}]
  wire [63:0] _GEN_15 = 5'hf == io_reorderBuffer_0_bits_destinationRegister ? io_reorderBuffer_0_bits_value :
    registers_15; // @[RegisterFile.scala 37:26 46:{46,46}]
  wire [63:0] _GEN_16 = 5'h10 == io_reorderBuffer_0_bits_destinationRegister ? io_reorderBuffer_0_bits_value :
    registers_16; // @[RegisterFile.scala 37:26 46:{46,46}]
  wire [63:0] _GEN_17 = 5'h11 == io_reorderBuffer_0_bits_destinationRegister ? io_reorderBuffer_0_bits_value :
    registers_17; // @[RegisterFile.scala 37:26 46:{46,46}]
  wire [63:0] _GEN_18 = 5'h12 == io_reorderBuffer_0_bits_destinationRegister ? io_reorderBuffer_0_bits_value :
    registers_18; // @[RegisterFile.scala 37:26 46:{46,46}]
  wire [63:0] _GEN_19 = 5'h13 == io_reorderBuffer_0_bits_destinationRegister ? io_reorderBuffer_0_bits_value :
    registers_19; // @[RegisterFile.scala 37:26 46:{46,46}]
  wire [63:0] _GEN_20 = 5'h14 == io_reorderBuffer_0_bits_destinationRegister ? io_reorderBuffer_0_bits_value :
    registers_20; // @[RegisterFile.scala 37:26 46:{46,46}]
  wire [63:0] _GEN_21 = 5'h15 == io_reorderBuffer_0_bits_destinationRegister ? io_reorderBuffer_0_bits_value :
    registers_21; // @[RegisterFile.scala 37:26 46:{46,46}]
  wire [63:0] _GEN_22 = 5'h16 == io_reorderBuffer_0_bits_destinationRegister ? io_reorderBuffer_0_bits_value :
    registers_22; // @[RegisterFile.scala 37:26 46:{46,46}]
  wire [63:0] _GEN_23 = 5'h17 == io_reorderBuffer_0_bits_destinationRegister ? io_reorderBuffer_0_bits_value :
    registers_23; // @[RegisterFile.scala 37:26 46:{46,46}]
  wire [63:0] _GEN_24 = 5'h18 == io_reorderBuffer_0_bits_destinationRegister ? io_reorderBuffer_0_bits_value :
    registers_24; // @[RegisterFile.scala 37:26 46:{46,46}]
  wire [63:0] _GEN_25 = 5'h19 == io_reorderBuffer_0_bits_destinationRegister ? io_reorderBuffer_0_bits_value :
    registers_25; // @[RegisterFile.scala 37:26 46:{46,46}]
  wire [63:0] _GEN_26 = 5'h1a == io_reorderBuffer_0_bits_destinationRegister ? io_reorderBuffer_0_bits_value :
    registers_26; // @[RegisterFile.scala 37:26 46:{46,46}]
  wire [63:0] _GEN_27 = 5'h1b == io_reorderBuffer_0_bits_destinationRegister ? io_reorderBuffer_0_bits_value :
    registers_27; // @[RegisterFile.scala 37:26 46:{46,46}]
  wire [63:0] _GEN_28 = 5'h1c == io_reorderBuffer_0_bits_destinationRegister ? io_reorderBuffer_0_bits_value :
    registers_28; // @[RegisterFile.scala 37:26 46:{46,46}]
  wire [63:0] _GEN_29 = 5'h1d == io_reorderBuffer_0_bits_destinationRegister ? io_reorderBuffer_0_bits_value :
    registers_29; // @[RegisterFile.scala 37:26 46:{46,46}]
  wire [63:0] _GEN_30 = 5'h1e == io_reorderBuffer_0_bits_destinationRegister ? io_reorderBuffer_0_bits_value :
    registers_30; // @[RegisterFile.scala 37:26 46:{46,46}]
  wire [63:0] _GEN_31 = 5'h1f == io_reorderBuffer_0_bits_destinationRegister ? io_reorderBuffer_0_bits_value :
    registers_31; // @[RegisterFile.scala 37:26 46:{46,46}]
  wire [63:0] _GEN_33 = io_reorderBuffer_0_valid ? _GEN_1 : registers_1; // @[RegisterFile.scala 45:20 37:26]
  wire [63:0] _GEN_34 = io_reorderBuffer_0_valid ? _GEN_2 : registers_2; // @[RegisterFile.scala 45:20 37:26]
  wire [63:0] _GEN_35 = io_reorderBuffer_0_valid ? _GEN_3 : registers_3; // @[RegisterFile.scala 45:20 37:26]
  wire [63:0] _GEN_36 = io_reorderBuffer_0_valid ? _GEN_4 : registers_4; // @[RegisterFile.scala 45:20 37:26]
  wire [63:0] _GEN_37 = io_reorderBuffer_0_valid ? _GEN_5 : registers_5; // @[RegisterFile.scala 45:20 37:26]
  wire [63:0] _GEN_38 = io_reorderBuffer_0_valid ? _GEN_6 : registers_6; // @[RegisterFile.scala 45:20 37:26]
  wire [63:0] _GEN_39 = io_reorderBuffer_0_valid ? _GEN_7 : registers_7; // @[RegisterFile.scala 45:20 37:26]
  wire [63:0] _GEN_40 = io_reorderBuffer_0_valid ? _GEN_8 : registers_8; // @[RegisterFile.scala 45:20 37:26]
  wire [63:0] _GEN_41 = io_reorderBuffer_0_valid ? _GEN_9 : registers_9; // @[RegisterFile.scala 45:20 37:26]
  wire [63:0] _GEN_42 = io_reorderBuffer_0_valid ? _GEN_10 : registers_10; // @[RegisterFile.scala 45:20 37:26]
  wire [63:0] _GEN_43 = io_reorderBuffer_0_valid ? _GEN_11 : registers_11; // @[RegisterFile.scala 45:20 37:26]
  wire [63:0] _GEN_44 = io_reorderBuffer_0_valid ? _GEN_12 : registers_12; // @[RegisterFile.scala 45:20 37:26]
  wire [63:0] _GEN_45 = io_reorderBuffer_0_valid ? _GEN_13 : registers_13; // @[RegisterFile.scala 45:20 37:26]
  wire [63:0] _GEN_46 = io_reorderBuffer_0_valid ? _GEN_14 : registers_14; // @[RegisterFile.scala 45:20 37:26]
  wire [63:0] _GEN_47 = io_reorderBuffer_0_valid ? _GEN_15 : registers_15; // @[RegisterFile.scala 45:20 37:26]
  wire [63:0] _GEN_48 = io_reorderBuffer_0_valid ? _GEN_16 : registers_16; // @[RegisterFile.scala 45:20 37:26]
  wire [63:0] _GEN_49 = io_reorderBuffer_0_valid ? _GEN_17 : registers_17; // @[RegisterFile.scala 45:20 37:26]
  wire [63:0] _GEN_50 = io_reorderBuffer_0_valid ? _GEN_18 : registers_18; // @[RegisterFile.scala 45:20 37:26]
  wire [63:0] _GEN_51 = io_reorderBuffer_0_valid ? _GEN_19 : registers_19; // @[RegisterFile.scala 45:20 37:26]
  wire [63:0] _GEN_52 = io_reorderBuffer_0_valid ? _GEN_20 : registers_20; // @[RegisterFile.scala 45:20 37:26]
  wire [63:0] _GEN_53 = io_reorderBuffer_0_valid ? _GEN_21 : registers_21; // @[RegisterFile.scala 45:20 37:26]
  wire [63:0] _GEN_54 = io_reorderBuffer_0_valid ? _GEN_22 : registers_22; // @[RegisterFile.scala 45:20 37:26]
  wire [63:0] _GEN_55 = io_reorderBuffer_0_valid ? _GEN_23 : registers_23; // @[RegisterFile.scala 45:20 37:26]
  wire [63:0] _GEN_56 = io_reorderBuffer_0_valid ? _GEN_24 : registers_24; // @[RegisterFile.scala 45:20 37:26]
  wire [63:0] _GEN_57 = io_reorderBuffer_0_valid ? _GEN_25 : registers_25; // @[RegisterFile.scala 45:20 37:26]
  wire [63:0] _GEN_58 = io_reorderBuffer_0_valid ? _GEN_26 : registers_26; // @[RegisterFile.scala 45:20 37:26]
  wire [63:0] _GEN_59 = io_reorderBuffer_0_valid ? _GEN_27 : registers_27; // @[RegisterFile.scala 45:20 37:26]
  wire [63:0] _GEN_60 = io_reorderBuffer_0_valid ? _GEN_28 : registers_28; // @[RegisterFile.scala 45:20 37:26]
  wire [63:0] _GEN_61 = io_reorderBuffer_0_valid ? _GEN_29 : registers_29; // @[RegisterFile.scala 45:20 37:26]
  wire [63:0] _GEN_62 = io_reorderBuffer_0_valid ? _GEN_30 : registers_30; // @[RegisterFile.scala 45:20 37:26]
  wire [63:0] _GEN_63 = io_reorderBuffer_0_valid ? _GEN_31 : registers_31; // @[RegisterFile.scala 45:20 37:26]
  wire [63:0] _GEN_65 = 5'h1 == io_reorderBuffer_1_bits_destinationRegister ? io_reorderBuffer_1_bits_value : _GEN_33; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_66 = 5'h2 == io_reorderBuffer_1_bits_destinationRegister ? io_reorderBuffer_1_bits_value : _GEN_34; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_67 = 5'h3 == io_reorderBuffer_1_bits_destinationRegister ? io_reorderBuffer_1_bits_value : _GEN_35; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_68 = 5'h4 == io_reorderBuffer_1_bits_destinationRegister ? io_reorderBuffer_1_bits_value : _GEN_36; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_69 = 5'h5 == io_reorderBuffer_1_bits_destinationRegister ? io_reorderBuffer_1_bits_value : _GEN_37; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_70 = 5'h6 == io_reorderBuffer_1_bits_destinationRegister ? io_reorderBuffer_1_bits_value : _GEN_38; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_71 = 5'h7 == io_reorderBuffer_1_bits_destinationRegister ? io_reorderBuffer_1_bits_value : _GEN_39; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_72 = 5'h8 == io_reorderBuffer_1_bits_destinationRegister ? io_reorderBuffer_1_bits_value : _GEN_40; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_73 = 5'h9 == io_reorderBuffer_1_bits_destinationRegister ? io_reorderBuffer_1_bits_value : _GEN_41; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_74 = 5'ha == io_reorderBuffer_1_bits_destinationRegister ? io_reorderBuffer_1_bits_value : _GEN_42; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_75 = 5'hb == io_reorderBuffer_1_bits_destinationRegister ? io_reorderBuffer_1_bits_value : _GEN_43; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_76 = 5'hc == io_reorderBuffer_1_bits_destinationRegister ? io_reorderBuffer_1_bits_value : _GEN_44; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_77 = 5'hd == io_reorderBuffer_1_bits_destinationRegister ? io_reorderBuffer_1_bits_value : _GEN_45; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_78 = 5'he == io_reorderBuffer_1_bits_destinationRegister ? io_reorderBuffer_1_bits_value : _GEN_46; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_79 = 5'hf == io_reorderBuffer_1_bits_destinationRegister ? io_reorderBuffer_1_bits_value : _GEN_47; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_80 = 5'h10 == io_reorderBuffer_1_bits_destinationRegister ? io_reorderBuffer_1_bits_value : _GEN_48; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_81 = 5'h11 == io_reorderBuffer_1_bits_destinationRegister ? io_reorderBuffer_1_bits_value : _GEN_49; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_82 = 5'h12 == io_reorderBuffer_1_bits_destinationRegister ? io_reorderBuffer_1_bits_value : _GEN_50; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_83 = 5'h13 == io_reorderBuffer_1_bits_destinationRegister ? io_reorderBuffer_1_bits_value : _GEN_51; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_84 = 5'h14 == io_reorderBuffer_1_bits_destinationRegister ? io_reorderBuffer_1_bits_value : _GEN_52; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_85 = 5'h15 == io_reorderBuffer_1_bits_destinationRegister ? io_reorderBuffer_1_bits_value : _GEN_53; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_86 = 5'h16 == io_reorderBuffer_1_bits_destinationRegister ? io_reorderBuffer_1_bits_value : _GEN_54; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_87 = 5'h17 == io_reorderBuffer_1_bits_destinationRegister ? io_reorderBuffer_1_bits_value : _GEN_55; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_88 = 5'h18 == io_reorderBuffer_1_bits_destinationRegister ? io_reorderBuffer_1_bits_value : _GEN_56; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_89 = 5'h19 == io_reorderBuffer_1_bits_destinationRegister ? io_reorderBuffer_1_bits_value : _GEN_57; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_90 = 5'h1a == io_reorderBuffer_1_bits_destinationRegister ? io_reorderBuffer_1_bits_value : _GEN_58; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_91 = 5'h1b == io_reorderBuffer_1_bits_destinationRegister ? io_reorderBuffer_1_bits_value : _GEN_59; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_92 = 5'h1c == io_reorderBuffer_1_bits_destinationRegister ? io_reorderBuffer_1_bits_value : _GEN_60; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_93 = 5'h1d == io_reorderBuffer_1_bits_destinationRegister ? io_reorderBuffer_1_bits_value : _GEN_61; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_94 = 5'h1e == io_reorderBuffer_1_bits_destinationRegister ? io_reorderBuffer_1_bits_value : _GEN_62; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_95 = 5'h1f == io_reorderBuffer_1_bits_destinationRegister ? io_reorderBuffer_1_bits_value : _GEN_63; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_97 = io_reorderBuffer_1_valid ? _GEN_65 : _GEN_33; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_98 = io_reorderBuffer_1_valid ? _GEN_66 : _GEN_34; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_99 = io_reorderBuffer_1_valid ? _GEN_67 : _GEN_35; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_100 = io_reorderBuffer_1_valid ? _GEN_68 : _GEN_36; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_101 = io_reorderBuffer_1_valid ? _GEN_69 : _GEN_37; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_102 = io_reorderBuffer_1_valid ? _GEN_70 : _GEN_38; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_103 = io_reorderBuffer_1_valid ? _GEN_71 : _GEN_39; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_104 = io_reorderBuffer_1_valid ? _GEN_72 : _GEN_40; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_105 = io_reorderBuffer_1_valid ? _GEN_73 : _GEN_41; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_106 = io_reorderBuffer_1_valid ? _GEN_74 : _GEN_42; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_107 = io_reorderBuffer_1_valid ? _GEN_75 : _GEN_43; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_108 = io_reorderBuffer_1_valid ? _GEN_76 : _GEN_44; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_109 = io_reorderBuffer_1_valid ? _GEN_77 : _GEN_45; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_110 = io_reorderBuffer_1_valid ? _GEN_78 : _GEN_46; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_111 = io_reorderBuffer_1_valid ? _GEN_79 : _GEN_47; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_112 = io_reorderBuffer_1_valid ? _GEN_80 : _GEN_48; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_113 = io_reorderBuffer_1_valid ? _GEN_81 : _GEN_49; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_114 = io_reorderBuffer_1_valid ? _GEN_82 : _GEN_50; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_115 = io_reorderBuffer_1_valid ? _GEN_83 : _GEN_51; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_116 = io_reorderBuffer_1_valid ? _GEN_84 : _GEN_52; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_117 = io_reorderBuffer_1_valid ? _GEN_85 : _GEN_53; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_118 = io_reorderBuffer_1_valid ? _GEN_86 : _GEN_54; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_119 = io_reorderBuffer_1_valid ? _GEN_87 : _GEN_55; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_120 = io_reorderBuffer_1_valid ? _GEN_88 : _GEN_56; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_121 = io_reorderBuffer_1_valid ? _GEN_89 : _GEN_57; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_122 = io_reorderBuffer_1_valid ? _GEN_90 : _GEN_58; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_123 = io_reorderBuffer_1_valid ? _GEN_91 : _GEN_59; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_124 = io_reorderBuffer_1_valid ? _GEN_92 : _GEN_60; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_125 = io_reorderBuffer_1_valid ? _GEN_93 : _GEN_61; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_126 = io_reorderBuffer_1_valid ? _GEN_94 : _GEN_62; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_127 = io_reorderBuffer_1_valid ? _GEN_95 : _GEN_63; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_129 = 5'h1 == io_reorderBuffer_2_bits_destinationRegister ? io_reorderBuffer_2_bits_value : _GEN_97; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_130 = 5'h2 == io_reorderBuffer_2_bits_destinationRegister ? io_reorderBuffer_2_bits_value : _GEN_98; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_131 = 5'h3 == io_reorderBuffer_2_bits_destinationRegister ? io_reorderBuffer_2_bits_value : _GEN_99; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_132 = 5'h4 == io_reorderBuffer_2_bits_destinationRegister ? io_reorderBuffer_2_bits_value : _GEN_100; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_133 = 5'h5 == io_reorderBuffer_2_bits_destinationRegister ? io_reorderBuffer_2_bits_value : _GEN_101; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_134 = 5'h6 == io_reorderBuffer_2_bits_destinationRegister ? io_reorderBuffer_2_bits_value : _GEN_102; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_135 = 5'h7 == io_reorderBuffer_2_bits_destinationRegister ? io_reorderBuffer_2_bits_value : _GEN_103; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_136 = 5'h8 == io_reorderBuffer_2_bits_destinationRegister ? io_reorderBuffer_2_bits_value : _GEN_104; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_137 = 5'h9 == io_reorderBuffer_2_bits_destinationRegister ? io_reorderBuffer_2_bits_value : _GEN_105; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_138 = 5'ha == io_reorderBuffer_2_bits_destinationRegister ? io_reorderBuffer_2_bits_value : _GEN_106; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_139 = 5'hb == io_reorderBuffer_2_bits_destinationRegister ? io_reorderBuffer_2_bits_value : _GEN_107; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_140 = 5'hc == io_reorderBuffer_2_bits_destinationRegister ? io_reorderBuffer_2_bits_value : _GEN_108; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_141 = 5'hd == io_reorderBuffer_2_bits_destinationRegister ? io_reorderBuffer_2_bits_value : _GEN_109; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_142 = 5'he == io_reorderBuffer_2_bits_destinationRegister ? io_reorderBuffer_2_bits_value : _GEN_110; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_143 = 5'hf == io_reorderBuffer_2_bits_destinationRegister ? io_reorderBuffer_2_bits_value : _GEN_111; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_144 = 5'h10 == io_reorderBuffer_2_bits_destinationRegister ? io_reorderBuffer_2_bits_value : _GEN_112
    ; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_145 = 5'h11 == io_reorderBuffer_2_bits_destinationRegister ? io_reorderBuffer_2_bits_value : _GEN_113
    ; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_146 = 5'h12 == io_reorderBuffer_2_bits_destinationRegister ? io_reorderBuffer_2_bits_value : _GEN_114
    ; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_147 = 5'h13 == io_reorderBuffer_2_bits_destinationRegister ? io_reorderBuffer_2_bits_value : _GEN_115
    ; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_148 = 5'h14 == io_reorderBuffer_2_bits_destinationRegister ? io_reorderBuffer_2_bits_value : _GEN_116
    ; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_149 = 5'h15 == io_reorderBuffer_2_bits_destinationRegister ? io_reorderBuffer_2_bits_value : _GEN_117
    ; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_150 = 5'h16 == io_reorderBuffer_2_bits_destinationRegister ? io_reorderBuffer_2_bits_value : _GEN_118
    ; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_151 = 5'h17 == io_reorderBuffer_2_bits_destinationRegister ? io_reorderBuffer_2_bits_value : _GEN_119
    ; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_152 = 5'h18 == io_reorderBuffer_2_bits_destinationRegister ? io_reorderBuffer_2_bits_value : _GEN_120
    ; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_153 = 5'h19 == io_reorderBuffer_2_bits_destinationRegister ? io_reorderBuffer_2_bits_value : _GEN_121
    ; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_154 = 5'h1a == io_reorderBuffer_2_bits_destinationRegister ? io_reorderBuffer_2_bits_value : _GEN_122
    ; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_155 = 5'h1b == io_reorderBuffer_2_bits_destinationRegister ? io_reorderBuffer_2_bits_value : _GEN_123
    ; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_156 = 5'h1c == io_reorderBuffer_2_bits_destinationRegister ? io_reorderBuffer_2_bits_value : _GEN_124
    ; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_157 = 5'h1d == io_reorderBuffer_2_bits_destinationRegister ? io_reorderBuffer_2_bits_value : _GEN_125
    ; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_158 = 5'h1e == io_reorderBuffer_2_bits_destinationRegister ? io_reorderBuffer_2_bits_value : _GEN_126
    ; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_159 = 5'h1f == io_reorderBuffer_2_bits_destinationRegister ? io_reorderBuffer_2_bits_value : _GEN_127
    ; // @[RegisterFile.scala 46:{46,46}]
  wire [63:0] _GEN_161 = io_reorderBuffer_2_valid ? _GEN_129 : _GEN_97; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_162 = io_reorderBuffer_2_valid ? _GEN_130 : _GEN_98; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_163 = io_reorderBuffer_2_valid ? _GEN_131 : _GEN_99; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_164 = io_reorderBuffer_2_valid ? _GEN_132 : _GEN_100; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_165 = io_reorderBuffer_2_valid ? _GEN_133 : _GEN_101; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_166 = io_reorderBuffer_2_valid ? _GEN_134 : _GEN_102; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_167 = io_reorderBuffer_2_valid ? _GEN_135 : _GEN_103; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_168 = io_reorderBuffer_2_valid ? _GEN_136 : _GEN_104; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_169 = io_reorderBuffer_2_valid ? _GEN_137 : _GEN_105; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_170 = io_reorderBuffer_2_valid ? _GEN_138 : _GEN_106; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_171 = io_reorderBuffer_2_valid ? _GEN_139 : _GEN_107; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_172 = io_reorderBuffer_2_valid ? _GEN_140 : _GEN_108; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_173 = io_reorderBuffer_2_valid ? _GEN_141 : _GEN_109; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_174 = io_reorderBuffer_2_valid ? _GEN_142 : _GEN_110; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_175 = io_reorderBuffer_2_valid ? _GEN_143 : _GEN_111; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_176 = io_reorderBuffer_2_valid ? _GEN_144 : _GEN_112; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_177 = io_reorderBuffer_2_valid ? _GEN_145 : _GEN_113; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_178 = io_reorderBuffer_2_valid ? _GEN_146 : _GEN_114; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_179 = io_reorderBuffer_2_valid ? _GEN_147 : _GEN_115; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_180 = io_reorderBuffer_2_valid ? _GEN_148 : _GEN_116; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_181 = io_reorderBuffer_2_valid ? _GEN_149 : _GEN_117; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_182 = io_reorderBuffer_2_valid ? _GEN_150 : _GEN_118; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_183 = io_reorderBuffer_2_valid ? _GEN_151 : _GEN_119; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_184 = io_reorderBuffer_2_valid ? _GEN_152 : _GEN_120; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_185 = io_reorderBuffer_2_valid ? _GEN_153 : _GEN_121; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_186 = io_reorderBuffer_2_valid ? _GEN_154 : _GEN_122; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_187 = io_reorderBuffer_2_valid ? _GEN_155 : _GEN_123; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_188 = io_reorderBuffer_2_valid ? _GEN_156 : _GEN_124; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_189 = io_reorderBuffer_2_valid ? _GEN_157 : _GEN_125; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_190 = io_reorderBuffer_2_valid ? _GEN_158 : _GEN_126; // @[RegisterFile.scala 45:20]
  wire [63:0] _GEN_191 = io_reorderBuffer_2_valid ? _GEN_159 : _GEN_127; // @[RegisterFile.scala 45:20]
  wire  _io_decoders_0_value1_T = io_decoders_0_sourceRegister1 == 5'h0; // @[RegisterFile.scala 54:27]
  wire [63:0] _GEN_257 = 5'h1 == io_decoders_0_sourceRegister1 ? registers_1 : 64'h0; // @[RegisterFile.scala 53:{22,22}]
  wire [63:0] _GEN_258 = 5'h2 == io_decoders_0_sourceRegister1 ? registers_2 : _GEN_257; // @[RegisterFile.scala 53:{22,22}]
  wire [63:0] _GEN_259 = 5'h3 == io_decoders_0_sourceRegister1 ? registers_3 : _GEN_258; // @[RegisterFile.scala 53:{22,22}]
  wire [63:0] _GEN_260 = 5'h4 == io_decoders_0_sourceRegister1 ? registers_4 : _GEN_259; // @[RegisterFile.scala 53:{22,22}]
  wire [63:0] _GEN_261 = 5'h5 == io_decoders_0_sourceRegister1 ? registers_5 : _GEN_260; // @[RegisterFile.scala 53:{22,22}]
  wire [63:0] _GEN_262 = 5'h6 == io_decoders_0_sourceRegister1 ? registers_6 : _GEN_261; // @[RegisterFile.scala 53:{22,22}]
  wire [63:0] _GEN_263 = 5'h7 == io_decoders_0_sourceRegister1 ? registers_7 : _GEN_262; // @[RegisterFile.scala 53:{22,22}]
  wire [63:0] _GEN_264 = 5'h8 == io_decoders_0_sourceRegister1 ? registers_8 : _GEN_263; // @[RegisterFile.scala 53:{22,22}]
  wire [63:0] _GEN_265 = 5'h9 == io_decoders_0_sourceRegister1 ? registers_9 : _GEN_264; // @[RegisterFile.scala 53:{22,22}]
  wire [63:0] _GEN_266 = 5'ha == io_decoders_0_sourceRegister1 ? registers_10 : _GEN_265; // @[RegisterFile.scala 53:{22,22}]
  wire [63:0] _GEN_267 = 5'hb == io_decoders_0_sourceRegister1 ? registers_11 : _GEN_266; // @[RegisterFile.scala 53:{22,22}]
  wire [63:0] _GEN_268 = 5'hc == io_decoders_0_sourceRegister1 ? registers_12 : _GEN_267; // @[RegisterFile.scala 53:{22,22}]
  wire [63:0] _GEN_269 = 5'hd == io_decoders_0_sourceRegister1 ? registers_13 : _GEN_268; // @[RegisterFile.scala 53:{22,22}]
  wire [63:0] _GEN_270 = 5'he == io_decoders_0_sourceRegister1 ? registers_14 : _GEN_269; // @[RegisterFile.scala 53:{22,22}]
  wire [63:0] _GEN_271 = 5'hf == io_decoders_0_sourceRegister1 ? registers_15 : _GEN_270; // @[RegisterFile.scala 53:{22,22}]
  wire [63:0] _GEN_272 = 5'h10 == io_decoders_0_sourceRegister1 ? registers_16 : _GEN_271; // @[RegisterFile.scala 53:{22,22}]
  wire [63:0] _GEN_273 = 5'h11 == io_decoders_0_sourceRegister1 ? registers_17 : _GEN_272; // @[RegisterFile.scala 53:{22,22}]
  wire [63:0] _GEN_274 = 5'h12 == io_decoders_0_sourceRegister1 ? registers_18 : _GEN_273; // @[RegisterFile.scala 53:{22,22}]
  wire [63:0] _GEN_275 = 5'h13 == io_decoders_0_sourceRegister1 ? registers_19 : _GEN_274; // @[RegisterFile.scala 53:{22,22}]
  wire [63:0] _GEN_276 = 5'h14 == io_decoders_0_sourceRegister1 ? registers_20 : _GEN_275; // @[RegisterFile.scala 53:{22,22}]
  wire [63:0] _GEN_277 = 5'h15 == io_decoders_0_sourceRegister1 ? registers_21 : _GEN_276; // @[RegisterFile.scala 53:{22,22}]
  wire [63:0] _GEN_278 = 5'h16 == io_decoders_0_sourceRegister1 ? registers_22 : _GEN_277; // @[RegisterFile.scala 53:{22,22}]
  wire [63:0] _GEN_279 = 5'h17 == io_decoders_0_sourceRegister1 ? registers_23 : _GEN_278; // @[RegisterFile.scala 53:{22,22}]
  wire [63:0] _GEN_280 = 5'h18 == io_decoders_0_sourceRegister1 ? registers_24 : _GEN_279; // @[RegisterFile.scala 53:{22,22}]
  wire [63:0] _GEN_281 = 5'h19 == io_decoders_0_sourceRegister1 ? registers_25 : _GEN_280; // @[RegisterFile.scala 53:{22,22}]
  wire [63:0] _GEN_282 = 5'h1a == io_decoders_0_sourceRegister1 ? registers_26 : _GEN_281; // @[RegisterFile.scala 53:{22,22}]
  wire [63:0] _GEN_283 = 5'h1b == io_decoders_0_sourceRegister1 ? registers_27 : _GEN_282; // @[RegisterFile.scala 53:{22,22}]
  wire [63:0] _GEN_284 = 5'h1c == io_decoders_0_sourceRegister1 ? registers_28 : _GEN_283; // @[RegisterFile.scala 53:{22,22}]
  wire [63:0] _GEN_285 = 5'h1d == io_decoders_0_sourceRegister1 ? registers_29 : _GEN_284; // @[RegisterFile.scala 53:{22,22}]
  wire [63:0] _GEN_286 = 5'h1e == io_decoders_0_sourceRegister1 ? registers_30 : _GEN_285; // @[RegisterFile.scala 53:{22,22}]
  wire [63:0] _GEN_287 = 5'h1f == io_decoders_0_sourceRegister1 ? registers_31 : _GEN_286; // @[RegisterFile.scala 53:{22,22}]
  wire  _io_decoders_0_value2_T = io_decoders_0_sourceRegister2 == 5'h0; // @[RegisterFile.scala 59:27]
  wire [63:0] _GEN_289 = 5'h1 == io_decoders_0_sourceRegister2 ? registers_1 : 64'h0; // @[RegisterFile.scala 58:{22,22}]
  wire [63:0] _GEN_290 = 5'h2 == io_decoders_0_sourceRegister2 ? registers_2 : _GEN_289; // @[RegisterFile.scala 58:{22,22}]
  wire [63:0] _GEN_291 = 5'h3 == io_decoders_0_sourceRegister2 ? registers_3 : _GEN_290; // @[RegisterFile.scala 58:{22,22}]
  wire [63:0] _GEN_292 = 5'h4 == io_decoders_0_sourceRegister2 ? registers_4 : _GEN_291; // @[RegisterFile.scala 58:{22,22}]
  wire [63:0] _GEN_293 = 5'h5 == io_decoders_0_sourceRegister2 ? registers_5 : _GEN_292; // @[RegisterFile.scala 58:{22,22}]
  wire [63:0] _GEN_294 = 5'h6 == io_decoders_0_sourceRegister2 ? registers_6 : _GEN_293; // @[RegisterFile.scala 58:{22,22}]
  wire [63:0] _GEN_295 = 5'h7 == io_decoders_0_sourceRegister2 ? registers_7 : _GEN_294; // @[RegisterFile.scala 58:{22,22}]
  wire [63:0] _GEN_296 = 5'h8 == io_decoders_0_sourceRegister2 ? registers_8 : _GEN_295; // @[RegisterFile.scala 58:{22,22}]
  wire [63:0] _GEN_297 = 5'h9 == io_decoders_0_sourceRegister2 ? registers_9 : _GEN_296; // @[RegisterFile.scala 58:{22,22}]
  wire [63:0] _GEN_298 = 5'ha == io_decoders_0_sourceRegister2 ? registers_10 : _GEN_297; // @[RegisterFile.scala 58:{22,22}]
  wire [63:0] _GEN_299 = 5'hb == io_decoders_0_sourceRegister2 ? registers_11 : _GEN_298; // @[RegisterFile.scala 58:{22,22}]
  wire [63:0] _GEN_300 = 5'hc == io_decoders_0_sourceRegister2 ? registers_12 : _GEN_299; // @[RegisterFile.scala 58:{22,22}]
  wire [63:0] _GEN_301 = 5'hd == io_decoders_0_sourceRegister2 ? registers_13 : _GEN_300; // @[RegisterFile.scala 58:{22,22}]
  wire [63:0] _GEN_302 = 5'he == io_decoders_0_sourceRegister2 ? registers_14 : _GEN_301; // @[RegisterFile.scala 58:{22,22}]
  wire [63:0] _GEN_303 = 5'hf == io_decoders_0_sourceRegister2 ? registers_15 : _GEN_302; // @[RegisterFile.scala 58:{22,22}]
  wire [63:0] _GEN_304 = 5'h10 == io_decoders_0_sourceRegister2 ? registers_16 : _GEN_303; // @[RegisterFile.scala 58:{22,22}]
  wire [63:0] _GEN_305 = 5'h11 == io_decoders_0_sourceRegister2 ? registers_17 : _GEN_304; // @[RegisterFile.scala 58:{22,22}]
  wire [63:0] _GEN_306 = 5'h12 == io_decoders_0_sourceRegister2 ? registers_18 : _GEN_305; // @[RegisterFile.scala 58:{22,22}]
  wire [63:0] _GEN_307 = 5'h13 == io_decoders_0_sourceRegister2 ? registers_19 : _GEN_306; // @[RegisterFile.scala 58:{22,22}]
  wire [63:0] _GEN_308 = 5'h14 == io_decoders_0_sourceRegister2 ? registers_20 : _GEN_307; // @[RegisterFile.scala 58:{22,22}]
  wire [63:0] _GEN_309 = 5'h15 == io_decoders_0_sourceRegister2 ? registers_21 : _GEN_308; // @[RegisterFile.scala 58:{22,22}]
  wire [63:0] _GEN_310 = 5'h16 == io_decoders_0_sourceRegister2 ? registers_22 : _GEN_309; // @[RegisterFile.scala 58:{22,22}]
  wire [63:0] _GEN_311 = 5'h17 == io_decoders_0_sourceRegister2 ? registers_23 : _GEN_310; // @[RegisterFile.scala 58:{22,22}]
  wire [63:0] _GEN_312 = 5'h18 == io_decoders_0_sourceRegister2 ? registers_24 : _GEN_311; // @[RegisterFile.scala 58:{22,22}]
  wire [63:0] _GEN_313 = 5'h19 == io_decoders_0_sourceRegister2 ? registers_25 : _GEN_312; // @[RegisterFile.scala 58:{22,22}]
  wire [63:0] _GEN_314 = 5'h1a == io_decoders_0_sourceRegister2 ? registers_26 : _GEN_313; // @[RegisterFile.scala 58:{22,22}]
  wire [63:0] _GEN_315 = 5'h1b == io_decoders_0_sourceRegister2 ? registers_27 : _GEN_314; // @[RegisterFile.scala 58:{22,22}]
  wire [63:0] _GEN_316 = 5'h1c == io_decoders_0_sourceRegister2 ? registers_28 : _GEN_315; // @[RegisterFile.scala 58:{22,22}]
  wire [63:0] _GEN_317 = 5'h1d == io_decoders_0_sourceRegister2 ? registers_29 : _GEN_316; // @[RegisterFile.scala 58:{22,22}]
  wire [63:0] _GEN_318 = 5'h1e == io_decoders_0_sourceRegister2 ? registers_30 : _GEN_317; // @[RegisterFile.scala 58:{22,22}]
  wire [63:0] _GEN_319 = 5'h1f == io_decoders_0_sourceRegister2 ? registers_31 : _GEN_318; // @[RegisterFile.scala 58:{22,22}]
  assign io_decoders_0_value1 = _io_decoders_0_value1_T ? 64'h0 : _GEN_287; // @[RegisterFile.scala 53:22]
  assign io_decoders_0_value2 = _io_decoders_0_value2_T ? 64'h0 : _GEN_319; // @[RegisterFile.scala 58:22]
  always @(posedge clock) begin
    if (reset) begin // @[RegisterFile.scala 37:26]
      registers_1 <= 64'h0; // @[RegisterFile.scala 37:26]
    end else if (io_reorderBuffer_3_valid) begin // @[RegisterFile.scala 45:20]
      if (5'h1 == io_reorderBuffer_3_bits_destinationRegister) begin // @[RegisterFile.scala 46:46]
        registers_1 <= io_reorderBuffer_3_bits_value; // @[RegisterFile.scala 46:46]
      end else begin
        registers_1 <= _GEN_161;
      end
    end else begin
      registers_1 <= _GEN_161;
    end
    if (reset) begin // @[RegisterFile.scala 37:26]
      registers_2 <= 64'h0; // @[RegisterFile.scala 37:26]
    end else if (io_reorderBuffer_3_valid) begin // @[RegisterFile.scala 45:20]
      if (5'h2 == io_reorderBuffer_3_bits_destinationRegister) begin // @[RegisterFile.scala 46:46]
        registers_2 <= io_reorderBuffer_3_bits_value; // @[RegisterFile.scala 46:46]
      end else begin
        registers_2 <= _GEN_162;
      end
    end else begin
      registers_2 <= _GEN_162;
    end
    if (reset) begin // @[RegisterFile.scala 37:26]
      registers_3 <= 64'h0; // @[RegisterFile.scala 37:26]
    end else if (io_reorderBuffer_3_valid) begin // @[RegisterFile.scala 45:20]
      if (5'h3 == io_reorderBuffer_3_bits_destinationRegister) begin // @[RegisterFile.scala 46:46]
        registers_3 <= io_reorderBuffer_3_bits_value; // @[RegisterFile.scala 46:46]
      end else begin
        registers_3 <= _GEN_163;
      end
    end else begin
      registers_3 <= _GEN_163;
    end
    if (reset) begin // @[RegisterFile.scala 37:26]
      registers_4 <= 64'h1; // @[RegisterFile.scala 37:26]
    end else if (io_reorderBuffer_3_valid) begin // @[RegisterFile.scala 45:20]
      if (5'h4 == io_reorderBuffer_3_bits_destinationRegister) begin // @[RegisterFile.scala 46:46]
        registers_4 <= io_reorderBuffer_3_bits_value; // @[RegisterFile.scala 46:46]
      end else begin
        registers_4 <= _GEN_164;
      end
    end else begin
      registers_4 <= _GEN_164;
    end
    if (reset) begin // @[RegisterFile.scala 37:26]
      registers_5 <= 64'h0; // @[RegisterFile.scala 37:26]
    end else if (io_reorderBuffer_3_valid) begin // @[RegisterFile.scala 45:20]
      if (5'h5 == io_reorderBuffer_3_bits_destinationRegister) begin // @[RegisterFile.scala 46:46]
        registers_5 <= io_reorderBuffer_3_bits_value; // @[RegisterFile.scala 46:46]
      end else begin
        registers_5 <= _GEN_165;
      end
    end else begin
      registers_5 <= _GEN_165;
    end
    if (reset) begin // @[RegisterFile.scala 37:26]
      registers_6 <= 64'h0; // @[RegisterFile.scala 37:26]
    end else if (io_reorderBuffer_3_valid) begin // @[RegisterFile.scala 45:20]
      if (5'h6 == io_reorderBuffer_3_bits_destinationRegister) begin // @[RegisterFile.scala 46:46]
        registers_6 <= io_reorderBuffer_3_bits_value; // @[RegisterFile.scala 46:46]
      end else begin
        registers_6 <= _GEN_166;
      end
    end else begin
      registers_6 <= _GEN_166;
    end
    if (reset) begin // @[RegisterFile.scala 37:26]
      registers_7 <= 64'h0; // @[RegisterFile.scala 37:26]
    end else if (io_reorderBuffer_3_valid) begin // @[RegisterFile.scala 45:20]
      if (5'h7 == io_reorderBuffer_3_bits_destinationRegister) begin // @[RegisterFile.scala 46:46]
        registers_7 <= io_reorderBuffer_3_bits_value; // @[RegisterFile.scala 46:46]
      end else begin
        registers_7 <= _GEN_167;
      end
    end else begin
      registers_7 <= _GEN_167;
    end
    if (reset) begin // @[RegisterFile.scala 37:26]
      registers_8 <= 64'h0; // @[RegisterFile.scala 37:26]
    end else if (io_reorderBuffer_3_valid) begin // @[RegisterFile.scala 45:20]
      if (5'h8 == io_reorderBuffer_3_bits_destinationRegister) begin // @[RegisterFile.scala 46:46]
        registers_8 <= io_reorderBuffer_3_bits_value; // @[RegisterFile.scala 46:46]
      end else begin
        registers_8 <= _GEN_168;
      end
    end else begin
      registers_8 <= _GEN_168;
    end
    if (reset) begin // @[RegisterFile.scala 37:26]
      registers_9 <= 64'h0; // @[RegisterFile.scala 37:26]
    end else if (io_reorderBuffer_3_valid) begin // @[RegisterFile.scala 45:20]
      if (5'h9 == io_reorderBuffer_3_bits_destinationRegister) begin // @[RegisterFile.scala 46:46]
        registers_9 <= io_reorderBuffer_3_bits_value; // @[RegisterFile.scala 46:46]
      end else begin
        registers_9 <= _GEN_169;
      end
    end else begin
      registers_9 <= _GEN_169;
    end
    if (reset) begin // @[RegisterFile.scala 37:26]
      registers_10 <= 64'h0; // @[RegisterFile.scala 37:26]
    end else if (io_reorderBuffer_3_valid) begin // @[RegisterFile.scala 45:20]
      if (5'ha == io_reorderBuffer_3_bits_destinationRegister) begin // @[RegisterFile.scala 46:46]
        registers_10 <= io_reorderBuffer_3_bits_value; // @[RegisterFile.scala 46:46]
      end else begin
        registers_10 <= _GEN_170;
      end
    end else begin
      registers_10 <= _GEN_170;
    end
    if (reset) begin // @[RegisterFile.scala 37:26]
      registers_11 <= 64'h0; // @[RegisterFile.scala 37:26]
    end else if (io_reorderBuffer_3_valid) begin // @[RegisterFile.scala 45:20]
      if (5'hb == io_reorderBuffer_3_bits_destinationRegister) begin // @[RegisterFile.scala 46:46]
        registers_11 <= io_reorderBuffer_3_bits_value; // @[RegisterFile.scala 46:46]
      end else begin
        registers_11 <= _GEN_171;
      end
    end else begin
      registers_11 <= _GEN_171;
    end
    if (reset) begin // @[RegisterFile.scala 37:26]
      registers_12 <= 64'h0; // @[RegisterFile.scala 37:26]
    end else if (io_reorderBuffer_3_valid) begin // @[RegisterFile.scala 45:20]
      if (5'hc == io_reorderBuffer_3_bits_destinationRegister) begin // @[RegisterFile.scala 46:46]
        registers_12 <= io_reorderBuffer_3_bits_value; // @[RegisterFile.scala 46:46]
      end else begin
        registers_12 <= _GEN_172;
      end
    end else begin
      registers_12 <= _GEN_172;
    end
    if (reset) begin // @[RegisterFile.scala 37:26]
      registers_13 <= 64'h0; // @[RegisterFile.scala 37:26]
    end else if (io_reorderBuffer_3_valid) begin // @[RegisterFile.scala 45:20]
      if (5'hd == io_reorderBuffer_3_bits_destinationRegister) begin // @[RegisterFile.scala 46:46]
        registers_13 <= io_reorderBuffer_3_bits_value; // @[RegisterFile.scala 46:46]
      end else begin
        registers_13 <= _GEN_173;
      end
    end else begin
      registers_13 <= _GEN_173;
    end
    if (reset) begin // @[RegisterFile.scala 37:26]
      registers_14 <= 64'h0; // @[RegisterFile.scala 37:26]
    end else if (io_reorderBuffer_3_valid) begin // @[RegisterFile.scala 45:20]
      if (5'he == io_reorderBuffer_3_bits_destinationRegister) begin // @[RegisterFile.scala 46:46]
        registers_14 <= io_reorderBuffer_3_bits_value; // @[RegisterFile.scala 46:46]
      end else begin
        registers_14 <= _GEN_174;
      end
    end else begin
      registers_14 <= _GEN_174;
    end
    if (reset) begin // @[RegisterFile.scala 37:26]
      registers_15 <= 64'h0; // @[RegisterFile.scala 37:26]
    end else if (io_reorderBuffer_3_valid) begin // @[RegisterFile.scala 45:20]
      if (5'hf == io_reorderBuffer_3_bits_destinationRegister) begin // @[RegisterFile.scala 46:46]
        registers_15 <= io_reorderBuffer_3_bits_value; // @[RegisterFile.scala 46:46]
      end else begin
        registers_15 <= _GEN_175;
      end
    end else begin
      registers_15 <= _GEN_175;
    end
    if (reset) begin // @[RegisterFile.scala 37:26]
      registers_16 <= 64'h0; // @[RegisterFile.scala 37:26]
    end else if (io_reorderBuffer_3_valid) begin // @[RegisterFile.scala 45:20]
      if (5'h10 == io_reorderBuffer_3_bits_destinationRegister) begin // @[RegisterFile.scala 46:46]
        registers_16 <= io_reorderBuffer_3_bits_value; // @[RegisterFile.scala 46:46]
      end else begin
        registers_16 <= _GEN_176;
      end
    end else begin
      registers_16 <= _GEN_176;
    end
    if (reset) begin // @[RegisterFile.scala 37:26]
      registers_17 <= 64'h0; // @[RegisterFile.scala 37:26]
    end else if (io_reorderBuffer_3_valid) begin // @[RegisterFile.scala 45:20]
      if (5'h11 == io_reorderBuffer_3_bits_destinationRegister) begin // @[RegisterFile.scala 46:46]
        registers_17 <= io_reorderBuffer_3_bits_value; // @[RegisterFile.scala 46:46]
      end else begin
        registers_17 <= _GEN_177;
      end
    end else begin
      registers_17 <= _GEN_177;
    end
    if (reset) begin // @[RegisterFile.scala 37:26]
      registers_18 <= 64'h0; // @[RegisterFile.scala 37:26]
    end else if (io_reorderBuffer_3_valid) begin // @[RegisterFile.scala 45:20]
      if (5'h12 == io_reorderBuffer_3_bits_destinationRegister) begin // @[RegisterFile.scala 46:46]
        registers_18 <= io_reorderBuffer_3_bits_value; // @[RegisterFile.scala 46:46]
      end else begin
        registers_18 <= _GEN_178;
      end
    end else begin
      registers_18 <= _GEN_178;
    end
    if (reset) begin // @[RegisterFile.scala 37:26]
      registers_19 <= 64'h0; // @[RegisterFile.scala 37:26]
    end else if (io_reorderBuffer_3_valid) begin // @[RegisterFile.scala 45:20]
      if (5'h13 == io_reorderBuffer_3_bits_destinationRegister) begin // @[RegisterFile.scala 46:46]
        registers_19 <= io_reorderBuffer_3_bits_value; // @[RegisterFile.scala 46:46]
      end else begin
        registers_19 <= _GEN_179;
      end
    end else begin
      registers_19 <= _GEN_179;
    end
    if (reset) begin // @[RegisterFile.scala 37:26]
      registers_20 <= 64'h0; // @[RegisterFile.scala 37:26]
    end else if (io_reorderBuffer_3_valid) begin // @[RegisterFile.scala 45:20]
      if (5'h14 == io_reorderBuffer_3_bits_destinationRegister) begin // @[RegisterFile.scala 46:46]
        registers_20 <= io_reorderBuffer_3_bits_value; // @[RegisterFile.scala 46:46]
      end else begin
        registers_20 <= _GEN_180;
      end
    end else begin
      registers_20 <= _GEN_180;
    end
    if (reset) begin // @[RegisterFile.scala 37:26]
      registers_21 <= 64'h0; // @[RegisterFile.scala 37:26]
    end else if (io_reorderBuffer_3_valid) begin // @[RegisterFile.scala 45:20]
      if (5'h15 == io_reorderBuffer_3_bits_destinationRegister) begin // @[RegisterFile.scala 46:46]
        registers_21 <= io_reorderBuffer_3_bits_value; // @[RegisterFile.scala 46:46]
      end else begin
        registers_21 <= _GEN_181;
      end
    end else begin
      registers_21 <= _GEN_181;
    end
    if (reset) begin // @[RegisterFile.scala 37:26]
      registers_22 <= 64'h0; // @[RegisterFile.scala 37:26]
    end else if (io_reorderBuffer_3_valid) begin // @[RegisterFile.scala 45:20]
      if (5'h16 == io_reorderBuffer_3_bits_destinationRegister) begin // @[RegisterFile.scala 46:46]
        registers_22 <= io_reorderBuffer_3_bits_value; // @[RegisterFile.scala 46:46]
      end else begin
        registers_22 <= _GEN_182;
      end
    end else begin
      registers_22 <= _GEN_182;
    end
    if (reset) begin // @[RegisterFile.scala 37:26]
      registers_23 <= 64'h0; // @[RegisterFile.scala 37:26]
    end else if (io_reorderBuffer_3_valid) begin // @[RegisterFile.scala 45:20]
      if (5'h17 == io_reorderBuffer_3_bits_destinationRegister) begin // @[RegisterFile.scala 46:46]
        registers_23 <= io_reorderBuffer_3_bits_value; // @[RegisterFile.scala 46:46]
      end else begin
        registers_23 <= _GEN_183;
      end
    end else begin
      registers_23 <= _GEN_183;
    end
    if (reset) begin // @[RegisterFile.scala 37:26]
      registers_24 <= 64'h0; // @[RegisterFile.scala 37:26]
    end else if (io_reorderBuffer_3_valid) begin // @[RegisterFile.scala 45:20]
      if (5'h18 == io_reorderBuffer_3_bits_destinationRegister) begin // @[RegisterFile.scala 46:46]
        registers_24 <= io_reorderBuffer_3_bits_value; // @[RegisterFile.scala 46:46]
      end else begin
        registers_24 <= _GEN_184;
      end
    end else begin
      registers_24 <= _GEN_184;
    end
    if (reset) begin // @[RegisterFile.scala 37:26]
      registers_25 <= 64'h0; // @[RegisterFile.scala 37:26]
    end else if (io_reorderBuffer_3_valid) begin // @[RegisterFile.scala 45:20]
      if (5'h19 == io_reorderBuffer_3_bits_destinationRegister) begin // @[RegisterFile.scala 46:46]
        registers_25 <= io_reorderBuffer_3_bits_value; // @[RegisterFile.scala 46:46]
      end else begin
        registers_25 <= _GEN_185;
      end
    end else begin
      registers_25 <= _GEN_185;
    end
    if (reset) begin // @[RegisterFile.scala 37:26]
      registers_26 <= 64'h0; // @[RegisterFile.scala 37:26]
    end else if (io_reorderBuffer_3_valid) begin // @[RegisterFile.scala 45:20]
      if (5'h1a == io_reorderBuffer_3_bits_destinationRegister) begin // @[RegisterFile.scala 46:46]
        registers_26 <= io_reorderBuffer_3_bits_value; // @[RegisterFile.scala 46:46]
      end else begin
        registers_26 <= _GEN_186;
      end
    end else begin
      registers_26 <= _GEN_186;
    end
    if (reset) begin // @[RegisterFile.scala 37:26]
      registers_27 <= 64'h0; // @[RegisterFile.scala 37:26]
    end else if (io_reorderBuffer_3_valid) begin // @[RegisterFile.scala 45:20]
      if (5'h1b == io_reorderBuffer_3_bits_destinationRegister) begin // @[RegisterFile.scala 46:46]
        registers_27 <= io_reorderBuffer_3_bits_value; // @[RegisterFile.scala 46:46]
      end else begin
        registers_27 <= _GEN_187;
      end
    end else begin
      registers_27 <= _GEN_187;
    end
    if (reset) begin // @[RegisterFile.scala 37:26]
      registers_28 <= 64'h0; // @[RegisterFile.scala 37:26]
    end else if (io_reorderBuffer_3_valid) begin // @[RegisterFile.scala 45:20]
      if (5'h1c == io_reorderBuffer_3_bits_destinationRegister) begin // @[RegisterFile.scala 46:46]
        registers_28 <= io_reorderBuffer_3_bits_value; // @[RegisterFile.scala 46:46]
      end else begin
        registers_28 <= _GEN_188;
      end
    end else begin
      registers_28 <= _GEN_188;
    end
    if (reset) begin // @[RegisterFile.scala 37:26]
      registers_29 <= 64'h0; // @[RegisterFile.scala 37:26]
    end else if (io_reorderBuffer_3_valid) begin // @[RegisterFile.scala 45:20]
      if (5'h1d == io_reorderBuffer_3_bits_destinationRegister) begin // @[RegisterFile.scala 46:46]
        registers_29 <= io_reorderBuffer_3_bits_value; // @[RegisterFile.scala 46:46]
      end else begin
        registers_29 <= _GEN_189;
      end
    end else begin
      registers_29 <= _GEN_189;
    end
    if (reset) begin // @[RegisterFile.scala 37:26]
      registers_30 <= 64'h0; // @[RegisterFile.scala 37:26]
    end else if (io_reorderBuffer_3_valid) begin // @[RegisterFile.scala 45:20]
      if (5'h1e == io_reorderBuffer_3_bits_destinationRegister) begin // @[RegisterFile.scala 46:46]
        registers_30 <= io_reorderBuffer_3_bits_value; // @[RegisterFile.scala 46:46]
      end else begin
        registers_30 <= _GEN_190;
      end
    end else begin
      registers_30 <= _GEN_190;
    end
    if (reset) begin // @[RegisterFile.scala 37:26]
      registers_31 <= 64'h0; // @[RegisterFile.scala 37:26]
    end else if (io_reorderBuffer_3_valid) begin // @[RegisterFile.scala 45:20]
      if (5'h1f == io_reorderBuffer_3_bits_destinationRegister) begin // @[RegisterFile.scala 46:46]
        registers_31 <= io_reorderBuffer_3_bits_value; // @[RegisterFile.scala 46:46]
      end else begin
        registers_31 <= _GEN_191;
      end
    end else begin
      registers_31 <= _GEN_191;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  registers_1 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  registers_2 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  registers_3 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  registers_4 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  registers_5 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  registers_6 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  registers_7 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  registers_8 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  registers_9 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  registers_10 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  registers_11 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  registers_12 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  registers_13 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  registers_14 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  registers_15 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  registers_16 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  registers_17 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  registers_18 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  registers_19 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  registers_20 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  registers_21 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  registers_22 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  registers_23 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  registers_24 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  registers_25 = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  registers_26 = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  registers_27 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  registers_28 = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  registers_29 = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  registers_30 = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  registers_31 = _RAND_30[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module LoadStoreQueue(
  input         clock,
  input         reset,
  output        io_decoders_0_ready,
  input         io_decoders_0_valid,
  input         io_decoders_0_bits_accessInfo_accessType,
  input         io_decoders_0_bits_accessInfo_signed,
  input  [1:0]  io_decoders_0_bits_accessInfo_accessWidth,
  input         io_decoders_0_bits_addressAndLoadResultTag_threadId,
  input  [3:0]  io_decoders_0_bits_addressAndLoadResultTag_id,
  input  [63:0] io_decoders_0_bits_address,
  input         io_decoders_0_bits_addressValid,
  input         io_decoders_0_bits_storeDataTag_threadId,
  input  [3:0]  io_decoders_0_bits_storeDataTag_id,
  input  [63:0] io_decoders_0_bits_storeData,
  input         io_decoders_0_bits_storeDataValid,
  input         io_outputCollector_outputs_valid,
  input         io_outputCollector_outputs_bits_resultType,
  input  [63:0] io_outputCollector_outputs_bits_value,
  input         io_outputCollector_outputs_bits_tag_threadId,
  input  [3:0]  io_outputCollector_outputs_bits_tag_id,
  input         io_reorderBuffer_0_valid,
  input         io_reorderBuffer_0_bits_destinationTag_threadId,
  input  [3:0]  io_reorderBuffer_0_bits_destinationTag_id,
  input         io_reorderBuffer_1_valid,
  input         io_reorderBuffer_1_bits_destinationTag_threadId,
  input  [3:0]  io_reorderBuffer_1_bits_destinationTag_id,
  input         io_reorderBuffer_2_valid,
  input         io_reorderBuffer_2_bits_destinationTag_threadId,
  input  [3:0]  io_reorderBuffer_2_bits_destinationTag_id,
  input         io_reorderBuffer_3_valid,
  input         io_reorderBuffer_3_bits_destinationTag_threadId,
  input  [3:0]  io_reorderBuffer_3_bits_destinationTag_id,
  input         io_memory_ready,
  output        io_memory_valid,
  output [63:0] io_memory_bits_address,
  output        io_memory_bits_tag_threadId,
  output [3:0]  io_memory_bits_tag_id,
  output [63:0] io_memory_bits_data,
  output        io_memory_bits_accessInfo_accessType,
  output        io_memory_bits_accessInfo_signed,
  output [1:0]  io_memory_bits_accessInfo_accessWidth,
  output        io_isEmpty
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [63:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [63:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [63:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [63:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [63:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [63:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [63:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [63:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [63:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [63:0] _RAND_104;
  reg [31:0] _RAND_105;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] head; // @[LoadStoreQueue.scala 47:21]
  reg [2:0] nextTail; // @[LoadStoreQueue.scala 48:21]
  reg  buffer_0_valid; // @[LoadStoreQueue.scala 51:23]
  reg  buffer_0_readyReorderSign; // @[LoadStoreQueue.scala 51:23]
  reg  buffer_0_info_accessType; // @[LoadStoreQueue.scala 51:23]
  reg  buffer_0_info_signed; // @[LoadStoreQueue.scala 51:23]
  reg [1:0] buffer_0_info_accessWidth; // @[LoadStoreQueue.scala 51:23]
  reg  buffer_0_addressAndLoadResultTag_threadId; // @[LoadStoreQueue.scala 51:23]
  reg [3:0] buffer_0_addressAndLoadResultTag_id; // @[LoadStoreQueue.scala 51:23]
  reg [63:0] buffer_0_address; // @[LoadStoreQueue.scala 51:23]
  reg  buffer_0_addressValid; // @[LoadStoreQueue.scala 51:23]
  reg  buffer_0_storeDataTag_threadId; // @[LoadStoreQueue.scala 51:23]
  reg [3:0] buffer_0_storeDataTag_id; // @[LoadStoreQueue.scala 51:23]
  reg [63:0] buffer_0_storeData; // @[LoadStoreQueue.scala 51:23]
  reg  buffer_0_storeDataValid; // @[LoadStoreQueue.scala 51:23]
  reg  buffer_1_valid; // @[LoadStoreQueue.scala 51:23]
  reg  buffer_1_readyReorderSign; // @[LoadStoreQueue.scala 51:23]
  reg  buffer_1_info_accessType; // @[LoadStoreQueue.scala 51:23]
  reg  buffer_1_info_signed; // @[LoadStoreQueue.scala 51:23]
  reg [1:0] buffer_1_info_accessWidth; // @[LoadStoreQueue.scala 51:23]
  reg  buffer_1_addressAndLoadResultTag_threadId; // @[LoadStoreQueue.scala 51:23]
  reg [3:0] buffer_1_addressAndLoadResultTag_id; // @[LoadStoreQueue.scala 51:23]
  reg [63:0] buffer_1_address; // @[LoadStoreQueue.scala 51:23]
  reg  buffer_1_addressValid; // @[LoadStoreQueue.scala 51:23]
  reg  buffer_1_storeDataTag_threadId; // @[LoadStoreQueue.scala 51:23]
  reg [3:0] buffer_1_storeDataTag_id; // @[LoadStoreQueue.scala 51:23]
  reg [63:0] buffer_1_storeData; // @[LoadStoreQueue.scala 51:23]
  reg  buffer_1_storeDataValid; // @[LoadStoreQueue.scala 51:23]
  reg  buffer_2_valid; // @[LoadStoreQueue.scala 51:23]
  reg  buffer_2_readyReorderSign; // @[LoadStoreQueue.scala 51:23]
  reg  buffer_2_info_accessType; // @[LoadStoreQueue.scala 51:23]
  reg  buffer_2_info_signed; // @[LoadStoreQueue.scala 51:23]
  reg [1:0] buffer_2_info_accessWidth; // @[LoadStoreQueue.scala 51:23]
  reg  buffer_2_addressAndLoadResultTag_threadId; // @[LoadStoreQueue.scala 51:23]
  reg [3:0] buffer_2_addressAndLoadResultTag_id; // @[LoadStoreQueue.scala 51:23]
  reg [63:0] buffer_2_address; // @[LoadStoreQueue.scala 51:23]
  reg  buffer_2_addressValid; // @[LoadStoreQueue.scala 51:23]
  reg  buffer_2_storeDataTag_threadId; // @[LoadStoreQueue.scala 51:23]
  reg [3:0] buffer_2_storeDataTag_id; // @[LoadStoreQueue.scala 51:23]
  reg [63:0] buffer_2_storeData; // @[LoadStoreQueue.scala 51:23]
  reg  buffer_2_storeDataValid; // @[LoadStoreQueue.scala 51:23]
  reg  buffer_3_valid; // @[LoadStoreQueue.scala 51:23]
  reg  buffer_3_readyReorderSign; // @[LoadStoreQueue.scala 51:23]
  reg  buffer_3_info_accessType; // @[LoadStoreQueue.scala 51:23]
  reg  buffer_3_info_signed; // @[LoadStoreQueue.scala 51:23]
  reg [1:0] buffer_3_info_accessWidth; // @[LoadStoreQueue.scala 51:23]
  reg  buffer_3_addressAndLoadResultTag_threadId; // @[LoadStoreQueue.scala 51:23]
  reg [3:0] buffer_3_addressAndLoadResultTag_id; // @[LoadStoreQueue.scala 51:23]
  reg [63:0] buffer_3_address; // @[LoadStoreQueue.scala 51:23]
  reg  buffer_3_addressValid; // @[LoadStoreQueue.scala 51:23]
  reg  buffer_3_storeDataTag_threadId; // @[LoadStoreQueue.scala 51:23]
  reg [3:0] buffer_3_storeDataTag_id; // @[LoadStoreQueue.scala 51:23]
  reg [63:0] buffer_3_storeData; // @[LoadStoreQueue.scala 51:23]
  reg  buffer_3_storeDataValid; // @[LoadStoreQueue.scala 51:23]
  reg  buffer_4_valid; // @[LoadStoreQueue.scala 51:23]
  reg  buffer_4_readyReorderSign; // @[LoadStoreQueue.scala 51:23]
  reg  buffer_4_info_accessType; // @[LoadStoreQueue.scala 51:23]
  reg  buffer_4_info_signed; // @[LoadStoreQueue.scala 51:23]
  reg [1:0] buffer_4_info_accessWidth; // @[LoadStoreQueue.scala 51:23]
  reg  buffer_4_addressAndLoadResultTag_threadId; // @[LoadStoreQueue.scala 51:23]
  reg [3:0] buffer_4_addressAndLoadResultTag_id; // @[LoadStoreQueue.scala 51:23]
  reg [63:0] buffer_4_address; // @[LoadStoreQueue.scala 51:23]
  reg  buffer_4_addressValid; // @[LoadStoreQueue.scala 51:23]
  reg  buffer_4_storeDataTag_threadId; // @[LoadStoreQueue.scala 51:23]
  reg [3:0] buffer_4_storeDataTag_id; // @[LoadStoreQueue.scala 51:23]
  reg [63:0] buffer_4_storeData; // @[LoadStoreQueue.scala 51:23]
  reg  buffer_4_storeDataValid; // @[LoadStoreQueue.scala 51:23]
  reg  buffer_5_valid; // @[LoadStoreQueue.scala 51:23]
  reg  buffer_5_readyReorderSign; // @[LoadStoreQueue.scala 51:23]
  reg  buffer_5_info_accessType; // @[LoadStoreQueue.scala 51:23]
  reg  buffer_5_info_signed; // @[LoadStoreQueue.scala 51:23]
  reg [1:0] buffer_5_info_accessWidth; // @[LoadStoreQueue.scala 51:23]
  reg  buffer_5_addressAndLoadResultTag_threadId; // @[LoadStoreQueue.scala 51:23]
  reg [3:0] buffer_5_addressAndLoadResultTag_id; // @[LoadStoreQueue.scala 51:23]
  reg [63:0] buffer_5_address; // @[LoadStoreQueue.scala 51:23]
  reg  buffer_5_addressValid; // @[LoadStoreQueue.scala 51:23]
  reg  buffer_5_storeDataTag_threadId; // @[LoadStoreQueue.scala 51:23]
  reg [3:0] buffer_5_storeDataTag_id; // @[LoadStoreQueue.scala 51:23]
  reg [63:0] buffer_5_storeData; // @[LoadStoreQueue.scala 51:23]
  reg  buffer_5_storeDataValid; // @[LoadStoreQueue.scala 51:23]
  reg  buffer_6_valid; // @[LoadStoreQueue.scala 51:23]
  reg  buffer_6_readyReorderSign; // @[LoadStoreQueue.scala 51:23]
  reg  buffer_6_info_accessType; // @[LoadStoreQueue.scala 51:23]
  reg  buffer_6_info_signed; // @[LoadStoreQueue.scala 51:23]
  reg [1:0] buffer_6_info_accessWidth; // @[LoadStoreQueue.scala 51:23]
  reg  buffer_6_addressAndLoadResultTag_threadId; // @[LoadStoreQueue.scala 51:23]
  reg [3:0] buffer_6_addressAndLoadResultTag_id; // @[LoadStoreQueue.scala 51:23]
  reg [63:0] buffer_6_address; // @[LoadStoreQueue.scala 51:23]
  reg  buffer_6_addressValid; // @[LoadStoreQueue.scala 51:23]
  reg  buffer_6_storeDataTag_threadId; // @[LoadStoreQueue.scala 51:23]
  reg [3:0] buffer_6_storeDataTag_id; // @[LoadStoreQueue.scala 51:23]
  reg [63:0] buffer_6_storeData; // @[LoadStoreQueue.scala 51:23]
  reg  buffer_6_storeDataValid; // @[LoadStoreQueue.scala 51:23]
  reg  buffer_7_valid; // @[LoadStoreQueue.scala 51:23]
  reg  buffer_7_readyReorderSign; // @[LoadStoreQueue.scala 51:23]
  reg  buffer_7_info_accessType; // @[LoadStoreQueue.scala 51:23]
  reg  buffer_7_info_signed; // @[LoadStoreQueue.scala 51:23]
  reg [1:0] buffer_7_info_accessWidth; // @[LoadStoreQueue.scala 51:23]
  reg  buffer_7_addressAndLoadResultTag_threadId; // @[LoadStoreQueue.scala 51:23]
  reg [3:0] buffer_7_addressAndLoadResultTag_id; // @[LoadStoreQueue.scala 51:23]
  reg [63:0] buffer_7_address; // @[LoadStoreQueue.scala 51:23]
  reg  buffer_7_addressValid; // @[LoadStoreQueue.scala 51:23]
  reg  buffer_7_storeDataTag_threadId; // @[LoadStoreQueue.scala 51:23]
  reg [3:0] buffer_7_storeDataTag_id; // @[LoadStoreQueue.scala 51:23]
  reg [63:0] buffer_7_storeData; // @[LoadStoreQueue.scala 51:23]
  reg  buffer_7_storeDataValid; // @[LoadStoreQueue.scala 51:23]
  wire [2:0] _io_decoders_0_ready_T_1 = head + 3'h1; // @[LoadStoreQueue.scala 61:43]
  wire  entryValid = io_decoders_0_ready & io_decoders_0_valid; // @[LoadStoreQueue.scala 62:36]
  wire  _GEN_0 = 3'h0 == head | buffer_0_valid; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire  _GEN_1 = 3'h1 == head | buffer_1_valid; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire  _GEN_2 = 3'h2 == head | buffer_2_valid; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire  _GEN_3 = 3'h3 == head | buffer_3_valid; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire  _GEN_4 = 3'h4 == head | buffer_4_valid; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire  _GEN_5 = 3'h5 == head | buffer_5_valid; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire  _GEN_6 = 3'h6 == head | buffer_6_valid; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire  _GEN_7 = 3'h7 == head | buffer_7_valid; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire  _GEN_8 = 3'h0 == head ? 1'h0 : buffer_0_readyReorderSign; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire  _GEN_9 = 3'h1 == head ? 1'h0 : buffer_1_readyReorderSign; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire  _GEN_10 = 3'h2 == head ? 1'h0 : buffer_2_readyReorderSign; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire  _GEN_11 = 3'h3 == head ? 1'h0 : buffer_3_readyReorderSign; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire  _GEN_12 = 3'h4 == head ? 1'h0 : buffer_4_readyReorderSign; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire  _GEN_13 = 3'h5 == head ? 1'h0 : buffer_5_readyReorderSign; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire  _GEN_14 = 3'h6 == head ? 1'h0 : buffer_6_readyReorderSign; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire  _GEN_15 = 3'h7 == head ? 1'h0 : buffer_7_readyReorderSign; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire  _GEN_16 = 3'h0 == head ? io_decoders_0_bits_accessInfo_accessType : buffer_0_info_accessType; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire  _GEN_17 = 3'h1 == head ? io_decoders_0_bits_accessInfo_accessType : buffer_1_info_accessType; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire  _GEN_18 = 3'h2 == head ? io_decoders_0_bits_accessInfo_accessType : buffer_2_info_accessType; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire  _GEN_19 = 3'h3 == head ? io_decoders_0_bits_accessInfo_accessType : buffer_3_info_accessType; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire  _GEN_20 = 3'h4 == head ? io_decoders_0_bits_accessInfo_accessType : buffer_4_info_accessType; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire  _GEN_21 = 3'h5 == head ? io_decoders_0_bits_accessInfo_accessType : buffer_5_info_accessType; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire  _GEN_22 = 3'h6 == head ? io_decoders_0_bits_accessInfo_accessType : buffer_6_info_accessType; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire  _GEN_23 = 3'h7 == head ? io_decoders_0_bits_accessInfo_accessType : buffer_7_info_accessType; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire  _GEN_24 = 3'h0 == head ? io_decoders_0_bits_accessInfo_signed : buffer_0_info_signed; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire  _GEN_25 = 3'h1 == head ? io_decoders_0_bits_accessInfo_signed : buffer_1_info_signed; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire  _GEN_26 = 3'h2 == head ? io_decoders_0_bits_accessInfo_signed : buffer_2_info_signed; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire  _GEN_27 = 3'h3 == head ? io_decoders_0_bits_accessInfo_signed : buffer_3_info_signed; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire  _GEN_28 = 3'h4 == head ? io_decoders_0_bits_accessInfo_signed : buffer_4_info_signed; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire  _GEN_29 = 3'h5 == head ? io_decoders_0_bits_accessInfo_signed : buffer_5_info_signed; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire  _GEN_30 = 3'h6 == head ? io_decoders_0_bits_accessInfo_signed : buffer_6_info_signed; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire  _GEN_31 = 3'h7 == head ? io_decoders_0_bits_accessInfo_signed : buffer_7_info_signed; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire [1:0] _GEN_32 = 3'h0 == head ? io_decoders_0_bits_accessInfo_accessWidth : buffer_0_info_accessWidth; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire [1:0] _GEN_33 = 3'h1 == head ? io_decoders_0_bits_accessInfo_accessWidth : buffer_1_info_accessWidth; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire [1:0] _GEN_34 = 3'h2 == head ? io_decoders_0_bits_accessInfo_accessWidth : buffer_2_info_accessWidth; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire [1:0] _GEN_35 = 3'h3 == head ? io_decoders_0_bits_accessInfo_accessWidth : buffer_3_info_accessWidth; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire [1:0] _GEN_36 = 3'h4 == head ? io_decoders_0_bits_accessInfo_accessWidth : buffer_4_info_accessWidth; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire [1:0] _GEN_37 = 3'h5 == head ? io_decoders_0_bits_accessInfo_accessWidth : buffer_5_info_accessWidth; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire [1:0] _GEN_38 = 3'h6 == head ? io_decoders_0_bits_accessInfo_accessWidth : buffer_6_info_accessWidth; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire [1:0] _GEN_39 = 3'h7 == head ? io_decoders_0_bits_accessInfo_accessWidth : buffer_7_info_accessWidth; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire  _GEN_40 = 3'h0 == head ? io_decoders_0_bits_addressAndLoadResultTag_threadId :
    buffer_0_addressAndLoadResultTag_threadId; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire  _GEN_41 = 3'h1 == head ? io_decoders_0_bits_addressAndLoadResultTag_threadId :
    buffer_1_addressAndLoadResultTag_threadId; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire  _GEN_42 = 3'h2 == head ? io_decoders_0_bits_addressAndLoadResultTag_threadId :
    buffer_2_addressAndLoadResultTag_threadId; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire  _GEN_43 = 3'h3 == head ? io_decoders_0_bits_addressAndLoadResultTag_threadId :
    buffer_3_addressAndLoadResultTag_threadId; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire  _GEN_44 = 3'h4 == head ? io_decoders_0_bits_addressAndLoadResultTag_threadId :
    buffer_4_addressAndLoadResultTag_threadId; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire  _GEN_45 = 3'h5 == head ? io_decoders_0_bits_addressAndLoadResultTag_threadId :
    buffer_5_addressAndLoadResultTag_threadId; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire  _GEN_46 = 3'h6 == head ? io_decoders_0_bits_addressAndLoadResultTag_threadId :
    buffer_6_addressAndLoadResultTag_threadId; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire  _GEN_47 = 3'h7 == head ? io_decoders_0_bits_addressAndLoadResultTag_threadId :
    buffer_7_addressAndLoadResultTag_threadId; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire [3:0] _GEN_48 = 3'h0 == head ? io_decoders_0_bits_addressAndLoadResultTag_id :
    buffer_0_addressAndLoadResultTag_id; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire [3:0] _GEN_49 = 3'h1 == head ? io_decoders_0_bits_addressAndLoadResultTag_id :
    buffer_1_addressAndLoadResultTag_id; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire [3:0] _GEN_50 = 3'h2 == head ? io_decoders_0_bits_addressAndLoadResultTag_id :
    buffer_2_addressAndLoadResultTag_id; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire [3:0] _GEN_51 = 3'h3 == head ? io_decoders_0_bits_addressAndLoadResultTag_id :
    buffer_3_addressAndLoadResultTag_id; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire [3:0] _GEN_52 = 3'h4 == head ? io_decoders_0_bits_addressAndLoadResultTag_id :
    buffer_4_addressAndLoadResultTag_id; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire [3:0] _GEN_53 = 3'h5 == head ? io_decoders_0_bits_addressAndLoadResultTag_id :
    buffer_5_addressAndLoadResultTag_id; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire [3:0] _GEN_54 = 3'h6 == head ? io_decoders_0_bits_addressAndLoadResultTag_id :
    buffer_6_addressAndLoadResultTag_id; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire [3:0] _GEN_55 = 3'h7 == head ? io_decoders_0_bits_addressAndLoadResultTag_id :
    buffer_7_addressAndLoadResultTag_id; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire [63:0] _GEN_56 = 3'h0 == head ? io_decoders_0_bits_address : buffer_0_address; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire [63:0] _GEN_57 = 3'h1 == head ? io_decoders_0_bits_address : buffer_1_address; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire [63:0] _GEN_58 = 3'h2 == head ? io_decoders_0_bits_address : buffer_2_address; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire [63:0] _GEN_59 = 3'h3 == head ? io_decoders_0_bits_address : buffer_3_address; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire [63:0] _GEN_60 = 3'h4 == head ? io_decoders_0_bits_address : buffer_4_address; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire [63:0] _GEN_61 = 3'h5 == head ? io_decoders_0_bits_address : buffer_5_address; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire [63:0] _GEN_62 = 3'h6 == head ? io_decoders_0_bits_address : buffer_6_address; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire [63:0] _GEN_63 = 3'h7 == head ? io_decoders_0_bits_address : buffer_7_address; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire  _GEN_64 = 3'h0 == head ? io_decoders_0_bits_addressValid : buffer_0_addressValid; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire  _GEN_65 = 3'h1 == head ? io_decoders_0_bits_addressValid : buffer_1_addressValid; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire  _GEN_66 = 3'h2 == head ? io_decoders_0_bits_addressValid : buffer_2_addressValid; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire  _GEN_67 = 3'h3 == head ? io_decoders_0_bits_addressValid : buffer_3_addressValid; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire  _GEN_68 = 3'h4 == head ? io_decoders_0_bits_addressValid : buffer_4_addressValid; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire  _GEN_69 = 3'h5 == head ? io_decoders_0_bits_addressValid : buffer_5_addressValid; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire  _GEN_70 = 3'h6 == head ? io_decoders_0_bits_addressValid : buffer_6_addressValid; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire  _GEN_71 = 3'h7 == head ? io_decoders_0_bits_addressValid : buffer_7_addressValid; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire  _GEN_72 = 3'h0 == head ? io_decoders_0_bits_storeDataTag_threadId : buffer_0_storeDataTag_threadId; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire  _GEN_73 = 3'h1 == head ? io_decoders_0_bits_storeDataTag_threadId : buffer_1_storeDataTag_threadId; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire  _GEN_74 = 3'h2 == head ? io_decoders_0_bits_storeDataTag_threadId : buffer_2_storeDataTag_threadId; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire  _GEN_75 = 3'h3 == head ? io_decoders_0_bits_storeDataTag_threadId : buffer_3_storeDataTag_threadId; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire  _GEN_76 = 3'h4 == head ? io_decoders_0_bits_storeDataTag_threadId : buffer_4_storeDataTag_threadId; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire  _GEN_77 = 3'h5 == head ? io_decoders_0_bits_storeDataTag_threadId : buffer_5_storeDataTag_threadId; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire  _GEN_78 = 3'h6 == head ? io_decoders_0_bits_storeDataTag_threadId : buffer_6_storeDataTag_threadId; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire  _GEN_79 = 3'h7 == head ? io_decoders_0_bits_storeDataTag_threadId : buffer_7_storeDataTag_threadId; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire [3:0] _GEN_80 = 3'h0 == head ? io_decoders_0_bits_storeDataTag_id : buffer_0_storeDataTag_id; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire [3:0] _GEN_81 = 3'h1 == head ? io_decoders_0_bits_storeDataTag_id : buffer_1_storeDataTag_id; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire [3:0] _GEN_82 = 3'h2 == head ? io_decoders_0_bits_storeDataTag_id : buffer_2_storeDataTag_id; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire [3:0] _GEN_83 = 3'h3 == head ? io_decoders_0_bits_storeDataTag_id : buffer_3_storeDataTag_id; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire [3:0] _GEN_84 = 3'h4 == head ? io_decoders_0_bits_storeDataTag_id : buffer_4_storeDataTag_id; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire [3:0] _GEN_85 = 3'h5 == head ? io_decoders_0_bits_storeDataTag_id : buffer_5_storeDataTag_id; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire [3:0] _GEN_86 = 3'h6 == head ? io_decoders_0_bits_storeDataTag_id : buffer_6_storeDataTag_id; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire [3:0] _GEN_87 = 3'h7 == head ? io_decoders_0_bits_storeDataTag_id : buffer_7_storeDataTag_id; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire [63:0] _GEN_88 = 3'h0 == head ? io_decoders_0_bits_storeData : buffer_0_storeData; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire [63:0] _GEN_89 = 3'h1 == head ? io_decoders_0_bits_storeData : buffer_1_storeData; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire [63:0] _GEN_90 = 3'h2 == head ? io_decoders_0_bits_storeData : buffer_2_storeData; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire [63:0] _GEN_91 = 3'h3 == head ? io_decoders_0_bits_storeData : buffer_3_storeData; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire [63:0] _GEN_92 = 3'h4 == head ? io_decoders_0_bits_storeData : buffer_4_storeData; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire [63:0] _GEN_93 = 3'h5 == head ? io_decoders_0_bits_storeData : buffer_5_storeData; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire [63:0] _GEN_94 = 3'h6 == head ? io_decoders_0_bits_storeData : buffer_6_storeData; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire [63:0] _GEN_95 = 3'h7 == head ? io_decoders_0_bits_storeData : buffer_7_storeData; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire  _GEN_96 = 3'h0 == head ? io_decoders_0_bits_storeDataValid : buffer_0_storeDataValid; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire  _GEN_97 = 3'h1 == head ? io_decoders_0_bits_storeDataValid : buffer_1_storeDataValid; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire  _GEN_98 = 3'h2 == head ? io_decoders_0_bits_storeDataValid : buffer_2_storeDataValid; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire  _GEN_99 = 3'h3 == head ? io_decoders_0_bits_storeDataValid : buffer_3_storeDataValid; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire  _GEN_100 = 3'h4 == head ? io_decoders_0_bits_storeDataValid : buffer_4_storeDataValid; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire  _GEN_101 = 3'h5 == head ? io_decoders_0_bits_storeDataValid : buffer_5_storeDataValid; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire  _GEN_102 = 3'h6 == head ? io_decoders_0_bits_storeDataValid : buffer_6_storeDataValid; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire  _GEN_103 = 3'h7 == head ? io_decoders_0_bits_storeDataValid : buffer_7_storeDataValid; // @[LoadStoreQueue.scala 51:23 70:{27,27}]
  wire  _GEN_104 = entryValid ? _GEN_0 : buffer_0_valid; // @[LoadStoreQueue.scala 68:22 51:23]
  wire  _GEN_105 = entryValid ? _GEN_1 : buffer_1_valid; // @[LoadStoreQueue.scala 68:22 51:23]
  wire  _GEN_106 = entryValid ? _GEN_2 : buffer_2_valid; // @[LoadStoreQueue.scala 68:22 51:23]
  wire  _GEN_107 = entryValid ? _GEN_3 : buffer_3_valid; // @[LoadStoreQueue.scala 68:22 51:23]
  wire  _GEN_108 = entryValid ? _GEN_4 : buffer_4_valid; // @[LoadStoreQueue.scala 68:22 51:23]
  wire  _GEN_109 = entryValid ? _GEN_5 : buffer_5_valid; // @[LoadStoreQueue.scala 68:22 51:23]
  wire  _GEN_110 = entryValid ? _GEN_6 : buffer_6_valid; // @[LoadStoreQueue.scala 68:22 51:23]
  wire  _GEN_111 = entryValid ? _GEN_7 : buffer_7_valid; // @[LoadStoreQueue.scala 68:22 51:23]
  wire  _GEN_112 = entryValid ? _GEN_8 : buffer_0_readyReorderSign; // @[LoadStoreQueue.scala 68:22 51:23]
  wire  _GEN_113 = entryValid ? _GEN_9 : buffer_1_readyReorderSign; // @[LoadStoreQueue.scala 68:22 51:23]
  wire  _GEN_114 = entryValid ? _GEN_10 : buffer_2_readyReorderSign; // @[LoadStoreQueue.scala 68:22 51:23]
  wire  _GEN_115 = entryValid ? _GEN_11 : buffer_3_readyReorderSign; // @[LoadStoreQueue.scala 68:22 51:23]
  wire  _GEN_116 = entryValid ? _GEN_12 : buffer_4_readyReorderSign; // @[LoadStoreQueue.scala 68:22 51:23]
  wire  _GEN_117 = entryValid ? _GEN_13 : buffer_5_readyReorderSign; // @[LoadStoreQueue.scala 68:22 51:23]
  wire  _GEN_118 = entryValid ? _GEN_14 : buffer_6_readyReorderSign; // @[LoadStoreQueue.scala 68:22 51:23]
  wire  _GEN_119 = entryValid ? _GEN_15 : buffer_7_readyReorderSign; // @[LoadStoreQueue.scala 68:22 51:23]
  wire  _GEN_120 = entryValid ? _GEN_16 : buffer_0_info_accessType; // @[LoadStoreQueue.scala 68:22 51:23]
  wire  _GEN_121 = entryValid ? _GEN_17 : buffer_1_info_accessType; // @[LoadStoreQueue.scala 68:22 51:23]
  wire  _GEN_122 = entryValid ? _GEN_18 : buffer_2_info_accessType; // @[LoadStoreQueue.scala 68:22 51:23]
  wire  _GEN_123 = entryValid ? _GEN_19 : buffer_3_info_accessType; // @[LoadStoreQueue.scala 68:22 51:23]
  wire  _GEN_124 = entryValid ? _GEN_20 : buffer_4_info_accessType; // @[LoadStoreQueue.scala 68:22 51:23]
  wire  _GEN_125 = entryValid ? _GEN_21 : buffer_5_info_accessType; // @[LoadStoreQueue.scala 68:22 51:23]
  wire  _GEN_126 = entryValid ? _GEN_22 : buffer_6_info_accessType; // @[LoadStoreQueue.scala 68:22 51:23]
  wire  _GEN_127 = entryValid ? _GEN_23 : buffer_7_info_accessType; // @[LoadStoreQueue.scala 68:22 51:23]
  wire  _GEN_128 = entryValid ? _GEN_24 : buffer_0_info_signed; // @[LoadStoreQueue.scala 68:22 51:23]
  wire  _GEN_129 = entryValid ? _GEN_25 : buffer_1_info_signed; // @[LoadStoreQueue.scala 68:22 51:23]
  wire  _GEN_130 = entryValid ? _GEN_26 : buffer_2_info_signed; // @[LoadStoreQueue.scala 68:22 51:23]
  wire  _GEN_131 = entryValid ? _GEN_27 : buffer_3_info_signed; // @[LoadStoreQueue.scala 68:22 51:23]
  wire  _GEN_132 = entryValid ? _GEN_28 : buffer_4_info_signed; // @[LoadStoreQueue.scala 68:22 51:23]
  wire  _GEN_133 = entryValid ? _GEN_29 : buffer_5_info_signed; // @[LoadStoreQueue.scala 68:22 51:23]
  wire  _GEN_134 = entryValid ? _GEN_30 : buffer_6_info_signed; // @[LoadStoreQueue.scala 68:22 51:23]
  wire  _GEN_135 = entryValid ? _GEN_31 : buffer_7_info_signed; // @[LoadStoreQueue.scala 68:22 51:23]
  wire [1:0] _GEN_136 = entryValid ? _GEN_32 : buffer_0_info_accessWidth; // @[LoadStoreQueue.scala 68:22 51:23]
  wire [1:0] _GEN_137 = entryValid ? _GEN_33 : buffer_1_info_accessWidth; // @[LoadStoreQueue.scala 68:22 51:23]
  wire [1:0] _GEN_138 = entryValid ? _GEN_34 : buffer_2_info_accessWidth; // @[LoadStoreQueue.scala 68:22 51:23]
  wire [1:0] _GEN_139 = entryValid ? _GEN_35 : buffer_3_info_accessWidth; // @[LoadStoreQueue.scala 68:22 51:23]
  wire [1:0] _GEN_140 = entryValid ? _GEN_36 : buffer_4_info_accessWidth; // @[LoadStoreQueue.scala 68:22 51:23]
  wire [1:0] _GEN_141 = entryValid ? _GEN_37 : buffer_5_info_accessWidth; // @[LoadStoreQueue.scala 68:22 51:23]
  wire [1:0] _GEN_142 = entryValid ? _GEN_38 : buffer_6_info_accessWidth; // @[LoadStoreQueue.scala 68:22 51:23]
  wire [1:0] _GEN_143 = entryValid ? _GEN_39 : buffer_7_info_accessWidth; // @[LoadStoreQueue.scala 68:22 51:23]
  wire  _GEN_144 = entryValid ? _GEN_40 : buffer_0_addressAndLoadResultTag_threadId; // @[LoadStoreQueue.scala 68:22 51:23]
  wire  _GEN_145 = entryValid ? _GEN_41 : buffer_1_addressAndLoadResultTag_threadId; // @[LoadStoreQueue.scala 68:22 51:23]
  wire  _GEN_146 = entryValid ? _GEN_42 : buffer_2_addressAndLoadResultTag_threadId; // @[LoadStoreQueue.scala 68:22 51:23]
  wire  _GEN_147 = entryValid ? _GEN_43 : buffer_3_addressAndLoadResultTag_threadId; // @[LoadStoreQueue.scala 68:22 51:23]
  wire  _GEN_148 = entryValid ? _GEN_44 : buffer_4_addressAndLoadResultTag_threadId; // @[LoadStoreQueue.scala 68:22 51:23]
  wire  _GEN_149 = entryValid ? _GEN_45 : buffer_5_addressAndLoadResultTag_threadId; // @[LoadStoreQueue.scala 68:22 51:23]
  wire  _GEN_150 = entryValid ? _GEN_46 : buffer_6_addressAndLoadResultTag_threadId; // @[LoadStoreQueue.scala 68:22 51:23]
  wire  _GEN_151 = entryValid ? _GEN_47 : buffer_7_addressAndLoadResultTag_threadId; // @[LoadStoreQueue.scala 68:22 51:23]
  wire [3:0] _GEN_152 = entryValid ? _GEN_48 : buffer_0_addressAndLoadResultTag_id; // @[LoadStoreQueue.scala 68:22 51:23]
  wire [3:0] _GEN_153 = entryValid ? _GEN_49 : buffer_1_addressAndLoadResultTag_id; // @[LoadStoreQueue.scala 68:22 51:23]
  wire [3:0] _GEN_154 = entryValid ? _GEN_50 : buffer_2_addressAndLoadResultTag_id; // @[LoadStoreQueue.scala 68:22 51:23]
  wire [3:0] _GEN_155 = entryValid ? _GEN_51 : buffer_3_addressAndLoadResultTag_id; // @[LoadStoreQueue.scala 68:22 51:23]
  wire [3:0] _GEN_156 = entryValid ? _GEN_52 : buffer_4_addressAndLoadResultTag_id; // @[LoadStoreQueue.scala 68:22 51:23]
  wire [3:0] _GEN_157 = entryValid ? _GEN_53 : buffer_5_addressAndLoadResultTag_id; // @[LoadStoreQueue.scala 68:22 51:23]
  wire [3:0] _GEN_158 = entryValid ? _GEN_54 : buffer_6_addressAndLoadResultTag_id; // @[LoadStoreQueue.scala 68:22 51:23]
  wire [3:0] _GEN_159 = entryValid ? _GEN_55 : buffer_7_addressAndLoadResultTag_id; // @[LoadStoreQueue.scala 68:22 51:23]
  wire [63:0] _GEN_160 = entryValid ? _GEN_56 : buffer_0_address; // @[LoadStoreQueue.scala 68:22 51:23]
  wire [63:0] _GEN_161 = entryValid ? _GEN_57 : buffer_1_address; // @[LoadStoreQueue.scala 68:22 51:23]
  wire [63:0] _GEN_162 = entryValid ? _GEN_58 : buffer_2_address; // @[LoadStoreQueue.scala 68:22 51:23]
  wire [63:0] _GEN_163 = entryValid ? _GEN_59 : buffer_3_address; // @[LoadStoreQueue.scala 68:22 51:23]
  wire [63:0] _GEN_164 = entryValid ? _GEN_60 : buffer_4_address; // @[LoadStoreQueue.scala 68:22 51:23]
  wire [63:0] _GEN_165 = entryValid ? _GEN_61 : buffer_5_address; // @[LoadStoreQueue.scala 68:22 51:23]
  wire [63:0] _GEN_166 = entryValid ? _GEN_62 : buffer_6_address; // @[LoadStoreQueue.scala 68:22 51:23]
  wire [63:0] _GEN_167 = entryValid ? _GEN_63 : buffer_7_address; // @[LoadStoreQueue.scala 68:22 51:23]
  wire  _GEN_168 = entryValid ? _GEN_64 : buffer_0_addressValid; // @[LoadStoreQueue.scala 68:22 51:23]
  wire  _GEN_169 = entryValid ? _GEN_65 : buffer_1_addressValid; // @[LoadStoreQueue.scala 68:22 51:23]
  wire  _GEN_170 = entryValid ? _GEN_66 : buffer_2_addressValid; // @[LoadStoreQueue.scala 68:22 51:23]
  wire  _GEN_171 = entryValid ? _GEN_67 : buffer_3_addressValid; // @[LoadStoreQueue.scala 68:22 51:23]
  wire  _GEN_172 = entryValid ? _GEN_68 : buffer_4_addressValid; // @[LoadStoreQueue.scala 68:22 51:23]
  wire  _GEN_173 = entryValid ? _GEN_69 : buffer_5_addressValid; // @[LoadStoreQueue.scala 68:22 51:23]
  wire  _GEN_174 = entryValid ? _GEN_70 : buffer_6_addressValid; // @[LoadStoreQueue.scala 68:22 51:23]
  wire  _GEN_175 = entryValid ? _GEN_71 : buffer_7_addressValid; // @[LoadStoreQueue.scala 68:22 51:23]
  wire  _GEN_176 = entryValid ? _GEN_72 : buffer_0_storeDataTag_threadId; // @[LoadStoreQueue.scala 68:22 51:23]
  wire  _GEN_177 = entryValid ? _GEN_73 : buffer_1_storeDataTag_threadId; // @[LoadStoreQueue.scala 68:22 51:23]
  wire  _GEN_178 = entryValid ? _GEN_74 : buffer_2_storeDataTag_threadId; // @[LoadStoreQueue.scala 68:22 51:23]
  wire  _GEN_179 = entryValid ? _GEN_75 : buffer_3_storeDataTag_threadId; // @[LoadStoreQueue.scala 68:22 51:23]
  wire  _GEN_180 = entryValid ? _GEN_76 : buffer_4_storeDataTag_threadId; // @[LoadStoreQueue.scala 68:22 51:23]
  wire  _GEN_181 = entryValid ? _GEN_77 : buffer_5_storeDataTag_threadId; // @[LoadStoreQueue.scala 68:22 51:23]
  wire  _GEN_182 = entryValid ? _GEN_78 : buffer_6_storeDataTag_threadId; // @[LoadStoreQueue.scala 68:22 51:23]
  wire  _GEN_183 = entryValid ? _GEN_79 : buffer_7_storeDataTag_threadId; // @[LoadStoreQueue.scala 68:22 51:23]
  wire [3:0] _GEN_184 = entryValid ? _GEN_80 : buffer_0_storeDataTag_id; // @[LoadStoreQueue.scala 68:22 51:23]
  wire [3:0] _GEN_185 = entryValid ? _GEN_81 : buffer_1_storeDataTag_id; // @[LoadStoreQueue.scala 68:22 51:23]
  wire [3:0] _GEN_186 = entryValid ? _GEN_82 : buffer_2_storeDataTag_id; // @[LoadStoreQueue.scala 68:22 51:23]
  wire [3:0] _GEN_187 = entryValid ? _GEN_83 : buffer_3_storeDataTag_id; // @[LoadStoreQueue.scala 68:22 51:23]
  wire [3:0] _GEN_188 = entryValid ? _GEN_84 : buffer_4_storeDataTag_id; // @[LoadStoreQueue.scala 68:22 51:23]
  wire [3:0] _GEN_189 = entryValid ? _GEN_85 : buffer_5_storeDataTag_id; // @[LoadStoreQueue.scala 68:22 51:23]
  wire [3:0] _GEN_190 = entryValid ? _GEN_86 : buffer_6_storeDataTag_id; // @[LoadStoreQueue.scala 68:22 51:23]
  wire [3:0] _GEN_191 = entryValid ? _GEN_87 : buffer_7_storeDataTag_id; // @[LoadStoreQueue.scala 68:22 51:23]
  wire [63:0] _GEN_192 = entryValid ? _GEN_88 : buffer_0_storeData; // @[LoadStoreQueue.scala 68:22 51:23]
  wire [63:0] _GEN_193 = entryValid ? _GEN_89 : buffer_1_storeData; // @[LoadStoreQueue.scala 68:22 51:23]
  wire [63:0] _GEN_194 = entryValid ? _GEN_90 : buffer_2_storeData; // @[LoadStoreQueue.scala 68:22 51:23]
  wire [63:0] _GEN_195 = entryValid ? _GEN_91 : buffer_3_storeData; // @[LoadStoreQueue.scala 68:22 51:23]
  wire [63:0] _GEN_196 = entryValid ? _GEN_92 : buffer_4_storeData; // @[LoadStoreQueue.scala 68:22 51:23]
  wire [63:0] _GEN_197 = entryValid ? _GEN_93 : buffer_5_storeData; // @[LoadStoreQueue.scala 68:22 51:23]
  wire [63:0] _GEN_198 = entryValid ? _GEN_94 : buffer_6_storeData; // @[LoadStoreQueue.scala 68:22 51:23]
  wire [63:0] _GEN_199 = entryValid ? _GEN_95 : buffer_7_storeData; // @[LoadStoreQueue.scala 68:22 51:23]
  wire  _GEN_200 = entryValid ? _GEN_96 : buffer_0_storeDataValid; // @[LoadStoreQueue.scala 68:22 51:23]
  wire  _GEN_201 = entryValid ? _GEN_97 : buffer_1_storeDataValid; // @[LoadStoreQueue.scala 68:22 51:23]
  wire  _GEN_202 = entryValid ? _GEN_98 : buffer_2_storeDataValid; // @[LoadStoreQueue.scala 68:22 51:23]
  wire  _GEN_203 = entryValid ? _GEN_99 : buffer_3_storeDataValid; // @[LoadStoreQueue.scala 68:22 51:23]
  wire  _GEN_204 = entryValid ? _GEN_100 : buffer_4_storeDataValid; // @[LoadStoreQueue.scala 68:22 51:23]
  wire  _GEN_205 = entryValid ? _GEN_101 : buffer_5_storeDataValid; // @[LoadStoreQueue.scala 68:22 51:23]
  wire  _GEN_206 = entryValid ? _GEN_102 : buffer_6_storeDataValid; // @[LoadStoreQueue.scala 68:22 51:23]
  wire  _GEN_207 = entryValid ? _GEN_103 : buffer_7_storeDataValid; // @[LoadStoreQueue.scala 68:22 51:23]
  wire [2:0] _GEN_1962 = {{2'd0}, entryValid}; // @[LoadStoreQueue.scala 81:31]
  wire [2:0] insertIndex = head + _GEN_1962; // @[LoadStoreQueue.scala 81:31]
  wire  _T_5 = buffer_0_addressAndLoadResultTag_id == io_outputCollector_outputs_bits_tag_id &
    buffer_0_addressAndLoadResultTag_threadId == io_outputCollector_outputs_bits_tag_threadId; // @[Tag.scala 13:25]
  wire  _T_7 = _T_5 & ~buffer_0_addressValid; // @[LoadStoreQueue.scala 93:59]
  wire [63:0] _GEN_208 = _T_7 ? io_outputCollector_outputs_bits_value : _GEN_160; // @[LoadStoreQueue.scala 94:11 95:23]
  wire  _GEN_209 = _T_7 | _GEN_168; // @[LoadStoreQueue.scala 94:11 96:28]
  wire [63:0] _GEN_210 = io_outputCollector_outputs_bits_resultType ? _GEN_208 : _GEN_160; // @[LoadStoreQueue.scala 91:68]
  wire  _GEN_211 = io_outputCollector_outputs_bits_resultType ? _GEN_209 : _GEN_168; // @[LoadStoreQueue.scala 91:68]
  wire  _T_11 = buffer_0_storeDataTag_id == io_outputCollector_outputs_bits_tag_id & buffer_0_storeDataTag_threadId ==
    io_outputCollector_outputs_bits_tag_threadId; // @[Tag.scala 13:25]
  wire [63:0] _GEN_212 = _T_11 & ~buffer_0_storeDataValid ? io_outputCollector_outputs_bits_value : _GEN_192; // @[LoadStoreQueue.scala 100:75 101:25]
  wire  _GEN_213 = _T_11 & ~buffer_0_storeDataValid | _GEN_200; // @[LoadStoreQueue.scala 100:75 102:30]
  wire [63:0] _GEN_214 = ~io_outputCollector_outputs_bits_resultType ? _GEN_212 : _GEN_192; // @[LoadStoreQueue.scala 99:58]
  wire  _GEN_215 = ~io_outputCollector_outputs_bits_resultType ? _GEN_213 : _GEN_200; // @[LoadStoreQueue.scala 99:58]
  wire [63:0] _GEN_216 = io_outputCollector_outputs_valid & buffer_0_valid ? _GEN_210 : _GEN_160; // @[LoadStoreQueue.scala 90:37]
  wire  _GEN_217 = io_outputCollector_outputs_valid & buffer_0_valid ? _GEN_211 : _GEN_168; // @[LoadStoreQueue.scala 90:37]
  wire [63:0] _GEN_218 = io_outputCollector_outputs_valid & buffer_0_valid ? _GEN_214 : _GEN_192; // @[LoadStoreQueue.scala 90:37]
  wire  _GEN_219 = io_outputCollector_outputs_valid & buffer_0_valid ? _GEN_215 : _GEN_200; // @[LoadStoreQueue.scala 90:37]
  wire  _T_18 = buffer_1_addressAndLoadResultTag_id == io_outputCollector_outputs_bits_tag_id &
    buffer_1_addressAndLoadResultTag_threadId == io_outputCollector_outputs_bits_tag_threadId; // @[Tag.scala 13:25]
  wire  _T_20 = _T_18 & ~buffer_1_addressValid; // @[LoadStoreQueue.scala 93:59]
  wire [63:0] _GEN_220 = _T_20 ? io_outputCollector_outputs_bits_value : _GEN_161; // @[LoadStoreQueue.scala 94:11 95:23]
  wire  _GEN_221 = _T_20 | _GEN_169; // @[LoadStoreQueue.scala 94:11 96:28]
  wire [63:0] _GEN_222 = io_outputCollector_outputs_bits_resultType ? _GEN_220 : _GEN_161; // @[LoadStoreQueue.scala 91:68]
  wire  _GEN_223 = io_outputCollector_outputs_bits_resultType ? _GEN_221 : _GEN_169; // @[LoadStoreQueue.scala 91:68]
  wire  _T_24 = buffer_1_storeDataTag_id == io_outputCollector_outputs_bits_tag_id & buffer_1_storeDataTag_threadId ==
    io_outputCollector_outputs_bits_tag_threadId; // @[Tag.scala 13:25]
  wire [63:0] _GEN_224 = _T_24 & ~buffer_1_storeDataValid ? io_outputCollector_outputs_bits_value : _GEN_193; // @[LoadStoreQueue.scala 100:75 101:25]
  wire  _GEN_225 = _T_24 & ~buffer_1_storeDataValid | _GEN_201; // @[LoadStoreQueue.scala 100:75 102:30]
  wire [63:0] _GEN_226 = ~io_outputCollector_outputs_bits_resultType ? _GEN_224 : _GEN_193; // @[LoadStoreQueue.scala 99:58]
  wire  _GEN_227 = ~io_outputCollector_outputs_bits_resultType ? _GEN_225 : _GEN_201; // @[LoadStoreQueue.scala 99:58]
  wire [63:0] _GEN_228 = io_outputCollector_outputs_valid & buffer_1_valid ? _GEN_222 : _GEN_161; // @[LoadStoreQueue.scala 90:37]
  wire  _GEN_229 = io_outputCollector_outputs_valid & buffer_1_valid ? _GEN_223 : _GEN_169; // @[LoadStoreQueue.scala 90:37]
  wire [63:0] _GEN_230 = io_outputCollector_outputs_valid & buffer_1_valid ? _GEN_226 : _GEN_193; // @[LoadStoreQueue.scala 90:37]
  wire  _GEN_231 = io_outputCollector_outputs_valid & buffer_1_valid ? _GEN_227 : _GEN_201; // @[LoadStoreQueue.scala 90:37]
  wire  _T_31 = buffer_2_addressAndLoadResultTag_id == io_outputCollector_outputs_bits_tag_id &
    buffer_2_addressAndLoadResultTag_threadId == io_outputCollector_outputs_bits_tag_threadId; // @[Tag.scala 13:25]
  wire  _T_33 = _T_31 & ~buffer_2_addressValid; // @[LoadStoreQueue.scala 93:59]
  wire [63:0] _GEN_232 = _T_33 ? io_outputCollector_outputs_bits_value : _GEN_162; // @[LoadStoreQueue.scala 94:11 95:23]
  wire  _GEN_233 = _T_33 | _GEN_170; // @[LoadStoreQueue.scala 94:11 96:28]
  wire [63:0] _GEN_234 = io_outputCollector_outputs_bits_resultType ? _GEN_232 : _GEN_162; // @[LoadStoreQueue.scala 91:68]
  wire  _GEN_235 = io_outputCollector_outputs_bits_resultType ? _GEN_233 : _GEN_170; // @[LoadStoreQueue.scala 91:68]
  wire  _T_37 = buffer_2_storeDataTag_id == io_outputCollector_outputs_bits_tag_id & buffer_2_storeDataTag_threadId ==
    io_outputCollector_outputs_bits_tag_threadId; // @[Tag.scala 13:25]
  wire [63:0] _GEN_236 = _T_37 & ~buffer_2_storeDataValid ? io_outputCollector_outputs_bits_value : _GEN_194; // @[LoadStoreQueue.scala 100:75 101:25]
  wire  _GEN_237 = _T_37 & ~buffer_2_storeDataValid | _GEN_202; // @[LoadStoreQueue.scala 100:75 102:30]
  wire [63:0] _GEN_238 = ~io_outputCollector_outputs_bits_resultType ? _GEN_236 : _GEN_194; // @[LoadStoreQueue.scala 99:58]
  wire  _GEN_239 = ~io_outputCollector_outputs_bits_resultType ? _GEN_237 : _GEN_202; // @[LoadStoreQueue.scala 99:58]
  wire [63:0] _GEN_240 = io_outputCollector_outputs_valid & buffer_2_valid ? _GEN_234 : _GEN_162; // @[LoadStoreQueue.scala 90:37]
  wire  _GEN_241 = io_outputCollector_outputs_valid & buffer_2_valid ? _GEN_235 : _GEN_170; // @[LoadStoreQueue.scala 90:37]
  wire [63:0] _GEN_242 = io_outputCollector_outputs_valid & buffer_2_valid ? _GEN_238 : _GEN_194; // @[LoadStoreQueue.scala 90:37]
  wire  _GEN_243 = io_outputCollector_outputs_valid & buffer_2_valid ? _GEN_239 : _GEN_202; // @[LoadStoreQueue.scala 90:37]
  wire  _T_44 = buffer_3_addressAndLoadResultTag_id == io_outputCollector_outputs_bits_tag_id &
    buffer_3_addressAndLoadResultTag_threadId == io_outputCollector_outputs_bits_tag_threadId; // @[Tag.scala 13:25]
  wire  _T_46 = _T_44 & ~buffer_3_addressValid; // @[LoadStoreQueue.scala 93:59]
  wire [63:0] _GEN_244 = _T_46 ? io_outputCollector_outputs_bits_value : _GEN_163; // @[LoadStoreQueue.scala 94:11 95:23]
  wire  _GEN_245 = _T_46 | _GEN_171; // @[LoadStoreQueue.scala 94:11 96:28]
  wire [63:0] _GEN_246 = io_outputCollector_outputs_bits_resultType ? _GEN_244 : _GEN_163; // @[LoadStoreQueue.scala 91:68]
  wire  _GEN_247 = io_outputCollector_outputs_bits_resultType ? _GEN_245 : _GEN_171; // @[LoadStoreQueue.scala 91:68]
  wire  _T_50 = buffer_3_storeDataTag_id == io_outputCollector_outputs_bits_tag_id & buffer_3_storeDataTag_threadId ==
    io_outputCollector_outputs_bits_tag_threadId; // @[Tag.scala 13:25]
  wire [63:0] _GEN_248 = _T_50 & ~buffer_3_storeDataValid ? io_outputCollector_outputs_bits_value : _GEN_195; // @[LoadStoreQueue.scala 100:75 101:25]
  wire  _GEN_249 = _T_50 & ~buffer_3_storeDataValid | _GEN_203; // @[LoadStoreQueue.scala 100:75 102:30]
  wire [63:0] _GEN_250 = ~io_outputCollector_outputs_bits_resultType ? _GEN_248 : _GEN_195; // @[LoadStoreQueue.scala 99:58]
  wire  _GEN_251 = ~io_outputCollector_outputs_bits_resultType ? _GEN_249 : _GEN_203; // @[LoadStoreQueue.scala 99:58]
  wire [63:0] _GEN_252 = io_outputCollector_outputs_valid & buffer_3_valid ? _GEN_246 : _GEN_163; // @[LoadStoreQueue.scala 90:37]
  wire  _GEN_253 = io_outputCollector_outputs_valid & buffer_3_valid ? _GEN_247 : _GEN_171; // @[LoadStoreQueue.scala 90:37]
  wire [63:0] _GEN_254 = io_outputCollector_outputs_valid & buffer_3_valid ? _GEN_250 : _GEN_195; // @[LoadStoreQueue.scala 90:37]
  wire  _GEN_255 = io_outputCollector_outputs_valid & buffer_3_valid ? _GEN_251 : _GEN_203; // @[LoadStoreQueue.scala 90:37]
  wire  _T_57 = buffer_4_addressAndLoadResultTag_id == io_outputCollector_outputs_bits_tag_id &
    buffer_4_addressAndLoadResultTag_threadId == io_outputCollector_outputs_bits_tag_threadId; // @[Tag.scala 13:25]
  wire  _T_59 = _T_57 & ~buffer_4_addressValid; // @[LoadStoreQueue.scala 93:59]
  wire [63:0] _GEN_256 = _T_59 ? io_outputCollector_outputs_bits_value : _GEN_164; // @[LoadStoreQueue.scala 94:11 95:23]
  wire  _GEN_257 = _T_59 | _GEN_172; // @[LoadStoreQueue.scala 94:11 96:28]
  wire [63:0] _GEN_258 = io_outputCollector_outputs_bits_resultType ? _GEN_256 : _GEN_164; // @[LoadStoreQueue.scala 91:68]
  wire  _GEN_259 = io_outputCollector_outputs_bits_resultType ? _GEN_257 : _GEN_172; // @[LoadStoreQueue.scala 91:68]
  wire  _T_63 = buffer_4_storeDataTag_id == io_outputCollector_outputs_bits_tag_id & buffer_4_storeDataTag_threadId ==
    io_outputCollector_outputs_bits_tag_threadId; // @[Tag.scala 13:25]
  wire [63:0] _GEN_260 = _T_63 & ~buffer_4_storeDataValid ? io_outputCollector_outputs_bits_value : _GEN_196; // @[LoadStoreQueue.scala 100:75 101:25]
  wire  _GEN_261 = _T_63 & ~buffer_4_storeDataValid | _GEN_204; // @[LoadStoreQueue.scala 100:75 102:30]
  wire [63:0] _GEN_262 = ~io_outputCollector_outputs_bits_resultType ? _GEN_260 : _GEN_196; // @[LoadStoreQueue.scala 99:58]
  wire  _GEN_263 = ~io_outputCollector_outputs_bits_resultType ? _GEN_261 : _GEN_204; // @[LoadStoreQueue.scala 99:58]
  wire [63:0] _GEN_264 = io_outputCollector_outputs_valid & buffer_4_valid ? _GEN_258 : _GEN_164; // @[LoadStoreQueue.scala 90:37]
  wire  _GEN_265 = io_outputCollector_outputs_valid & buffer_4_valid ? _GEN_259 : _GEN_172; // @[LoadStoreQueue.scala 90:37]
  wire [63:0] _GEN_266 = io_outputCollector_outputs_valid & buffer_4_valid ? _GEN_262 : _GEN_196; // @[LoadStoreQueue.scala 90:37]
  wire  _GEN_267 = io_outputCollector_outputs_valid & buffer_4_valid ? _GEN_263 : _GEN_204; // @[LoadStoreQueue.scala 90:37]
  wire  _T_70 = buffer_5_addressAndLoadResultTag_id == io_outputCollector_outputs_bits_tag_id &
    buffer_5_addressAndLoadResultTag_threadId == io_outputCollector_outputs_bits_tag_threadId; // @[Tag.scala 13:25]
  wire  _T_72 = _T_70 & ~buffer_5_addressValid; // @[LoadStoreQueue.scala 93:59]
  wire [63:0] _GEN_268 = _T_72 ? io_outputCollector_outputs_bits_value : _GEN_165; // @[LoadStoreQueue.scala 94:11 95:23]
  wire  _GEN_269 = _T_72 | _GEN_173; // @[LoadStoreQueue.scala 94:11 96:28]
  wire [63:0] _GEN_270 = io_outputCollector_outputs_bits_resultType ? _GEN_268 : _GEN_165; // @[LoadStoreQueue.scala 91:68]
  wire  _GEN_271 = io_outputCollector_outputs_bits_resultType ? _GEN_269 : _GEN_173; // @[LoadStoreQueue.scala 91:68]
  wire  _T_76 = buffer_5_storeDataTag_id == io_outputCollector_outputs_bits_tag_id & buffer_5_storeDataTag_threadId ==
    io_outputCollector_outputs_bits_tag_threadId; // @[Tag.scala 13:25]
  wire [63:0] _GEN_272 = _T_76 & ~buffer_5_storeDataValid ? io_outputCollector_outputs_bits_value : _GEN_197; // @[LoadStoreQueue.scala 100:75 101:25]
  wire  _GEN_273 = _T_76 & ~buffer_5_storeDataValid | _GEN_205; // @[LoadStoreQueue.scala 100:75 102:30]
  wire [63:0] _GEN_274 = ~io_outputCollector_outputs_bits_resultType ? _GEN_272 : _GEN_197; // @[LoadStoreQueue.scala 99:58]
  wire  _GEN_275 = ~io_outputCollector_outputs_bits_resultType ? _GEN_273 : _GEN_205; // @[LoadStoreQueue.scala 99:58]
  wire [63:0] _GEN_276 = io_outputCollector_outputs_valid & buffer_5_valid ? _GEN_270 : _GEN_165; // @[LoadStoreQueue.scala 90:37]
  wire  _GEN_277 = io_outputCollector_outputs_valid & buffer_5_valid ? _GEN_271 : _GEN_173; // @[LoadStoreQueue.scala 90:37]
  wire [63:0] _GEN_278 = io_outputCollector_outputs_valid & buffer_5_valid ? _GEN_274 : _GEN_197; // @[LoadStoreQueue.scala 90:37]
  wire  _GEN_279 = io_outputCollector_outputs_valid & buffer_5_valid ? _GEN_275 : _GEN_205; // @[LoadStoreQueue.scala 90:37]
  wire  _T_83 = buffer_6_addressAndLoadResultTag_id == io_outputCollector_outputs_bits_tag_id &
    buffer_6_addressAndLoadResultTag_threadId == io_outputCollector_outputs_bits_tag_threadId; // @[Tag.scala 13:25]
  wire  _T_85 = _T_83 & ~buffer_6_addressValid; // @[LoadStoreQueue.scala 93:59]
  wire [63:0] _GEN_280 = _T_85 ? io_outputCollector_outputs_bits_value : _GEN_166; // @[LoadStoreQueue.scala 94:11 95:23]
  wire  _GEN_281 = _T_85 | _GEN_174; // @[LoadStoreQueue.scala 94:11 96:28]
  wire [63:0] _GEN_282 = io_outputCollector_outputs_bits_resultType ? _GEN_280 : _GEN_166; // @[LoadStoreQueue.scala 91:68]
  wire  _GEN_283 = io_outputCollector_outputs_bits_resultType ? _GEN_281 : _GEN_174; // @[LoadStoreQueue.scala 91:68]
  wire  _T_89 = buffer_6_storeDataTag_id == io_outputCollector_outputs_bits_tag_id & buffer_6_storeDataTag_threadId ==
    io_outputCollector_outputs_bits_tag_threadId; // @[Tag.scala 13:25]
  wire [63:0] _GEN_284 = _T_89 & ~buffer_6_storeDataValid ? io_outputCollector_outputs_bits_value : _GEN_198; // @[LoadStoreQueue.scala 100:75 101:25]
  wire  _GEN_285 = _T_89 & ~buffer_6_storeDataValid | _GEN_206; // @[LoadStoreQueue.scala 100:75 102:30]
  wire [63:0] _GEN_286 = ~io_outputCollector_outputs_bits_resultType ? _GEN_284 : _GEN_198; // @[LoadStoreQueue.scala 99:58]
  wire  _GEN_287 = ~io_outputCollector_outputs_bits_resultType ? _GEN_285 : _GEN_206; // @[LoadStoreQueue.scala 99:58]
  wire [63:0] _GEN_288 = io_outputCollector_outputs_valid & buffer_6_valid ? _GEN_282 : _GEN_166; // @[LoadStoreQueue.scala 90:37]
  wire  _GEN_289 = io_outputCollector_outputs_valid & buffer_6_valid ? _GEN_283 : _GEN_174; // @[LoadStoreQueue.scala 90:37]
  wire [63:0] _GEN_290 = io_outputCollector_outputs_valid & buffer_6_valid ? _GEN_286 : _GEN_198; // @[LoadStoreQueue.scala 90:37]
  wire  _GEN_291 = io_outputCollector_outputs_valid & buffer_6_valid ? _GEN_287 : _GEN_206; // @[LoadStoreQueue.scala 90:37]
  wire  _T_96 = buffer_7_addressAndLoadResultTag_id == io_outputCollector_outputs_bits_tag_id &
    buffer_7_addressAndLoadResultTag_threadId == io_outputCollector_outputs_bits_tag_threadId; // @[Tag.scala 13:25]
  wire  _T_98 = _T_96 & ~buffer_7_addressValid; // @[LoadStoreQueue.scala 93:59]
  wire [63:0] _GEN_292 = _T_98 ? io_outputCollector_outputs_bits_value : _GEN_167; // @[LoadStoreQueue.scala 94:11 95:23]
  wire  _GEN_293 = _T_98 | _GEN_175; // @[LoadStoreQueue.scala 94:11 96:28]
  wire [63:0] _GEN_294 = io_outputCollector_outputs_bits_resultType ? _GEN_292 : _GEN_167; // @[LoadStoreQueue.scala 91:68]
  wire  _GEN_295 = io_outputCollector_outputs_bits_resultType ? _GEN_293 : _GEN_175; // @[LoadStoreQueue.scala 91:68]
  wire  _T_102 = buffer_7_storeDataTag_id == io_outputCollector_outputs_bits_tag_id & buffer_7_storeDataTag_threadId ==
    io_outputCollector_outputs_bits_tag_threadId; // @[Tag.scala 13:25]
  wire [63:0] _GEN_296 = _T_102 & ~buffer_7_storeDataValid ? io_outputCollector_outputs_bits_value : _GEN_199; // @[LoadStoreQueue.scala 100:75 101:25]
  wire  _GEN_297 = _T_102 & ~buffer_7_storeDataValid | _GEN_207; // @[LoadStoreQueue.scala 100:75 102:30]
  wire [63:0] _GEN_298 = ~io_outputCollector_outputs_bits_resultType ? _GEN_296 : _GEN_199; // @[LoadStoreQueue.scala 99:58]
  wire  _GEN_299 = ~io_outputCollector_outputs_bits_resultType ? _GEN_297 : _GEN_207; // @[LoadStoreQueue.scala 99:58]
  wire [63:0] _GEN_300 = io_outputCollector_outputs_valid & buffer_7_valid ? _GEN_294 : _GEN_167; // @[LoadStoreQueue.scala 90:37]
  wire  _GEN_301 = io_outputCollector_outputs_valid & buffer_7_valid ? _GEN_295 : _GEN_175; // @[LoadStoreQueue.scala 90:37]
  wire [63:0] _GEN_302 = io_outputCollector_outputs_valid & buffer_7_valid ? _GEN_298 : _GEN_199; // @[LoadStoreQueue.scala 90:37]
  wire  _GEN_303 = io_outputCollector_outputs_valid & buffer_7_valid ? _GEN_299 : _GEN_207; // @[LoadStoreQueue.scala 90:37]
  wire  _T_107 = io_reorderBuffer_0_bits_destinationTag_id == buffer_0_addressAndLoadResultTag_id &
    io_reorderBuffer_0_bits_destinationTag_threadId == buffer_0_addressAndLoadResultTag_threadId; // @[Tag.scala 13:25]
  wire  _T_108 = buffer_0_valid & _T_107; // @[LoadStoreQueue.scala 112:21]
  wire  _GEN_304 = _T_108 | _GEN_112; // @[LoadStoreQueue.scala 113:11 114:32]
  wire  _T_111 = io_reorderBuffer_0_bits_destinationTag_id == buffer_1_addressAndLoadResultTag_id &
    io_reorderBuffer_0_bits_destinationTag_threadId == buffer_1_addressAndLoadResultTag_threadId; // @[Tag.scala 13:25]
  wire  _T_112 = buffer_1_valid & _T_111; // @[LoadStoreQueue.scala 112:21]
  wire  _GEN_305 = _T_112 | _GEN_113; // @[LoadStoreQueue.scala 113:11 114:32]
  wire  _T_115 = io_reorderBuffer_0_bits_destinationTag_id == buffer_2_addressAndLoadResultTag_id &
    io_reorderBuffer_0_bits_destinationTag_threadId == buffer_2_addressAndLoadResultTag_threadId; // @[Tag.scala 13:25]
  wire  _T_116 = buffer_2_valid & _T_115; // @[LoadStoreQueue.scala 112:21]
  wire  _GEN_306 = _T_116 | _GEN_114; // @[LoadStoreQueue.scala 113:11 114:32]
  wire  _T_119 = io_reorderBuffer_0_bits_destinationTag_id == buffer_3_addressAndLoadResultTag_id &
    io_reorderBuffer_0_bits_destinationTag_threadId == buffer_3_addressAndLoadResultTag_threadId; // @[Tag.scala 13:25]
  wire  _T_120 = buffer_3_valid & _T_119; // @[LoadStoreQueue.scala 112:21]
  wire  _GEN_307 = _T_120 | _GEN_115; // @[LoadStoreQueue.scala 113:11 114:32]
  wire  _T_123 = io_reorderBuffer_0_bits_destinationTag_id == buffer_4_addressAndLoadResultTag_id &
    io_reorderBuffer_0_bits_destinationTag_threadId == buffer_4_addressAndLoadResultTag_threadId; // @[Tag.scala 13:25]
  wire  _T_124 = buffer_4_valid & _T_123; // @[LoadStoreQueue.scala 112:21]
  wire  _GEN_308 = _T_124 | _GEN_116; // @[LoadStoreQueue.scala 113:11 114:32]
  wire  _T_127 = io_reorderBuffer_0_bits_destinationTag_id == buffer_5_addressAndLoadResultTag_id &
    io_reorderBuffer_0_bits_destinationTag_threadId == buffer_5_addressAndLoadResultTag_threadId; // @[Tag.scala 13:25]
  wire  _T_128 = buffer_5_valid & _T_127; // @[LoadStoreQueue.scala 112:21]
  wire  _GEN_309 = _T_128 | _GEN_117; // @[LoadStoreQueue.scala 113:11 114:32]
  wire  _T_131 = io_reorderBuffer_0_bits_destinationTag_id == buffer_6_addressAndLoadResultTag_id &
    io_reorderBuffer_0_bits_destinationTag_threadId == buffer_6_addressAndLoadResultTag_threadId; // @[Tag.scala 13:25]
  wire  _T_132 = buffer_6_valid & _T_131; // @[LoadStoreQueue.scala 112:21]
  wire  _GEN_310 = _T_132 | _GEN_118; // @[LoadStoreQueue.scala 113:11 114:32]
  wire  _T_135 = io_reorderBuffer_0_bits_destinationTag_id == buffer_7_addressAndLoadResultTag_id &
    io_reorderBuffer_0_bits_destinationTag_threadId == buffer_7_addressAndLoadResultTag_threadId; // @[Tag.scala 13:25]
  wire  _T_136 = buffer_7_valid & _T_135; // @[LoadStoreQueue.scala 112:21]
  wire  _GEN_311 = _T_136 | _GEN_119; // @[LoadStoreQueue.scala 113:11 114:32]
  wire  _GEN_312 = io_reorderBuffer_0_valid ? _GEN_304 : _GEN_112; // @[LoadStoreQueue.scala 109:20]
  wire  _GEN_313 = io_reorderBuffer_0_valid ? _GEN_305 : _GEN_113; // @[LoadStoreQueue.scala 109:20]
  wire  _GEN_314 = io_reorderBuffer_0_valid ? _GEN_306 : _GEN_114; // @[LoadStoreQueue.scala 109:20]
  wire  _GEN_315 = io_reorderBuffer_0_valid ? _GEN_307 : _GEN_115; // @[LoadStoreQueue.scala 109:20]
  wire  _GEN_316 = io_reorderBuffer_0_valid ? _GEN_308 : _GEN_116; // @[LoadStoreQueue.scala 109:20]
  wire  _GEN_317 = io_reorderBuffer_0_valid ? _GEN_309 : _GEN_117; // @[LoadStoreQueue.scala 109:20]
  wire  _GEN_318 = io_reorderBuffer_0_valid ? _GEN_310 : _GEN_118; // @[LoadStoreQueue.scala 109:20]
  wire  _GEN_319 = io_reorderBuffer_0_valid ? _GEN_311 : _GEN_119; // @[LoadStoreQueue.scala 109:20]
  wire  _T_139 = io_reorderBuffer_1_bits_destinationTag_id == buffer_0_addressAndLoadResultTag_id &
    io_reorderBuffer_1_bits_destinationTag_threadId == buffer_0_addressAndLoadResultTag_threadId; // @[Tag.scala 13:25]
  wire  _T_140 = buffer_0_valid & _T_139; // @[LoadStoreQueue.scala 112:21]
  wire  _GEN_320 = _T_140 | _GEN_312; // @[LoadStoreQueue.scala 113:11 114:32]
  wire  _T_143 = io_reorderBuffer_1_bits_destinationTag_id == buffer_1_addressAndLoadResultTag_id &
    io_reorderBuffer_1_bits_destinationTag_threadId == buffer_1_addressAndLoadResultTag_threadId; // @[Tag.scala 13:25]
  wire  _T_144 = buffer_1_valid & _T_143; // @[LoadStoreQueue.scala 112:21]
  wire  _GEN_321 = _T_144 | _GEN_313; // @[LoadStoreQueue.scala 113:11 114:32]
  wire  _T_147 = io_reorderBuffer_1_bits_destinationTag_id == buffer_2_addressAndLoadResultTag_id &
    io_reorderBuffer_1_bits_destinationTag_threadId == buffer_2_addressAndLoadResultTag_threadId; // @[Tag.scala 13:25]
  wire  _T_148 = buffer_2_valid & _T_147; // @[LoadStoreQueue.scala 112:21]
  wire  _GEN_322 = _T_148 | _GEN_314; // @[LoadStoreQueue.scala 113:11 114:32]
  wire  _T_151 = io_reorderBuffer_1_bits_destinationTag_id == buffer_3_addressAndLoadResultTag_id &
    io_reorderBuffer_1_bits_destinationTag_threadId == buffer_3_addressAndLoadResultTag_threadId; // @[Tag.scala 13:25]
  wire  _T_152 = buffer_3_valid & _T_151; // @[LoadStoreQueue.scala 112:21]
  wire  _GEN_323 = _T_152 | _GEN_315; // @[LoadStoreQueue.scala 113:11 114:32]
  wire  _T_155 = io_reorderBuffer_1_bits_destinationTag_id == buffer_4_addressAndLoadResultTag_id &
    io_reorderBuffer_1_bits_destinationTag_threadId == buffer_4_addressAndLoadResultTag_threadId; // @[Tag.scala 13:25]
  wire  _T_156 = buffer_4_valid & _T_155; // @[LoadStoreQueue.scala 112:21]
  wire  _GEN_324 = _T_156 | _GEN_316; // @[LoadStoreQueue.scala 113:11 114:32]
  wire  _T_159 = io_reorderBuffer_1_bits_destinationTag_id == buffer_5_addressAndLoadResultTag_id &
    io_reorderBuffer_1_bits_destinationTag_threadId == buffer_5_addressAndLoadResultTag_threadId; // @[Tag.scala 13:25]
  wire  _T_160 = buffer_5_valid & _T_159; // @[LoadStoreQueue.scala 112:21]
  wire  _GEN_325 = _T_160 | _GEN_317; // @[LoadStoreQueue.scala 113:11 114:32]
  wire  _T_163 = io_reorderBuffer_1_bits_destinationTag_id == buffer_6_addressAndLoadResultTag_id &
    io_reorderBuffer_1_bits_destinationTag_threadId == buffer_6_addressAndLoadResultTag_threadId; // @[Tag.scala 13:25]
  wire  _T_164 = buffer_6_valid & _T_163; // @[LoadStoreQueue.scala 112:21]
  wire  _GEN_326 = _T_164 | _GEN_318; // @[LoadStoreQueue.scala 113:11 114:32]
  wire  _T_167 = io_reorderBuffer_1_bits_destinationTag_id == buffer_7_addressAndLoadResultTag_id &
    io_reorderBuffer_1_bits_destinationTag_threadId == buffer_7_addressAndLoadResultTag_threadId; // @[Tag.scala 13:25]
  wire  _T_168 = buffer_7_valid & _T_167; // @[LoadStoreQueue.scala 112:21]
  wire  _GEN_327 = _T_168 | _GEN_319; // @[LoadStoreQueue.scala 113:11 114:32]
  wire  _GEN_328 = io_reorderBuffer_1_valid ? _GEN_320 : _GEN_312; // @[LoadStoreQueue.scala 109:20]
  wire  _GEN_329 = io_reorderBuffer_1_valid ? _GEN_321 : _GEN_313; // @[LoadStoreQueue.scala 109:20]
  wire  _GEN_330 = io_reorderBuffer_1_valid ? _GEN_322 : _GEN_314; // @[LoadStoreQueue.scala 109:20]
  wire  _GEN_331 = io_reorderBuffer_1_valid ? _GEN_323 : _GEN_315; // @[LoadStoreQueue.scala 109:20]
  wire  _GEN_332 = io_reorderBuffer_1_valid ? _GEN_324 : _GEN_316; // @[LoadStoreQueue.scala 109:20]
  wire  _GEN_333 = io_reorderBuffer_1_valid ? _GEN_325 : _GEN_317; // @[LoadStoreQueue.scala 109:20]
  wire  _GEN_334 = io_reorderBuffer_1_valid ? _GEN_326 : _GEN_318; // @[LoadStoreQueue.scala 109:20]
  wire  _GEN_335 = io_reorderBuffer_1_valid ? _GEN_327 : _GEN_319; // @[LoadStoreQueue.scala 109:20]
  wire  _T_171 = io_reorderBuffer_2_bits_destinationTag_id == buffer_0_addressAndLoadResultTag_id &
    io_reorderBuffer_2_bits_destinationTag_threadId == buffer_0_addressAndLoadResultTag_threadId; // @[Tag.scala 13:25]
  wire  _T_172 = buffer_0_valid & _T_171; // @[LoadStoreQueue.scala 112:21]
  wire  _GEN_336 = _T_172 | _GEN_328; // @[LoadStoreQueue.scala 113:11 114:32]
  wire  _T_175 = io_reorderBuffer_2_bits_destinationTag_id == buffer_1_addressAndLoadResultTag_id &
    io_reorderBuffer_2_bits_destinationTag_threadId == buffer_1_addressAndLoadResultTag_threadId; // @[Tag.scala 13:25]
  wire  _T_176 = buffer_1_valid & _T_175; // @[LoadStoreQueue.scala 112:21]
  wire  _GEN_337 = _T_176 | _GEN_329; // @[LoadStoreQueue.scala 113:11 114:32]
  wire  _T_179 = io_reorderBuffer_2_bits_destinationTag_id == buffer_2_addressAndLoadResultTag_id &
    io_reorderBuffer_2_bits_destinationTag_threadId == buffer_2_addressAndLoadResultTag_threadId; // @[Tag.scala 13:25]
  wire  _T_180 = buffer_2_valid & _T_179; // @[LoadStoreQueue.scala 112:21]
  wire  _GEN_338 = _T_180 | _GEN_330; // @[LoadStoreQueue.scala 113:11 114:32]
  wire  _T_183 = io_reorderBuffer_2_bits_destinationTag_id == buffer_3_addressAndLoadResultTag_id &
    io_reorderBuffer_2_bits_destinationTag_threadId == buffer_3_addressAndLoadResultTag_threadId; // @[Tag.scala 13:25]
  wire  _T_184 = buffer_3_valid & _T_183; // @[LoadStoreQueue.scala 112:21]
  wire  _GEN_339 = _T_184 | _GEN_331; // @[LoadStoreQueue.scala 113:11 114:32]
  wire  _T_187 = io_reorderBuffer_2_bits_destinationTag_id == buffer_4_addressAndLoadResultTag_id &
    io_reorderBuffer_2_bits_destinationTag_threadId == buffer_4_addressAndLoadResultTag_threadId; // @[Tag.scala 13:25]
  wire  _T_188 = buffer_4_valid & _T_187; // @[LoadStoreQueue.scala 112:21]
  wire  _GEN_340 = _T_188 | _GEN_332; // @[LoadStoreQueue.scala 113:11 114:32]
  wire  _T_191 = io_reorderBuffer_2_bits_destinationTag_id == buffer_5_addressAndLoadResultTag_id &
    io_reorderBuffer_2_bits_destinationTag_threadId == buffer_5_addressAndLoadResultTag_threadId; // @[Tag.scala 13:25]
  wire  _T_192 = buffer_5_valid & _T_191; // @[LoadStoreQueue.scala 112:21]
  wire  _GEN_341 = _T_192 | _GEN_333; // @[LoadStoreQueue.scala 113:11 114:32]
  wire  _T_195 = io_reorderBuffer_2_bits_destinationTag_id == buffer_6_addressAndLoadResultTag_id &
    io_reorderBuffer_2_bits_destinationTag_threadId == buffer_6_addressAndLoadResultTag_threadId; // @[Tag.scala 13:25]
  wire  _T_196 = buffer_6_valid & _T_195; // @[LoadStoreQueue.scala 112:21]
  wire  _GEN_342 = _T_196 | _GEN_334; // @[LoadStoreQueue.scala 113:11 114:32]
  wire  _T_199 = io_reorderBuffer_2_bits_destinationTag_id == buffer_7_addressAndLoadResultTag_id &
    io_reorderBuffer_2_bits_destinationTag_threadId == buffer_7_addressAndLoadResultTag_threadId; // @[Tag.scala 13:25]
  wire  _T_200 = buffer_7_valid & _T_199; // @[LoadStoreQueue.scala 112:21]
  wire  _GEN_343 = _T_200 | _GEN_335; // @[LoadStoreQueue.scala 113:11 114:32]
  wire  _GEN_344 = io_reorderBuffer_2_valid ? _GEN_336 : _GEN_328; // @[LoadStoreQueue.scala 109:20]
  wire  _GEN_345 = io_reorderBuffer_2_valid ? _GEN_337 : _GEN_329; // @[LoadStoreQueue.scala 109:20]
  wire  _GEN_346 = io_reorderBuffer_2_valid ? _GEN_338 : _GEN_330; // @[LoadStoreQueue.scala 109:20]
  wire  _GEN_347 = io_reorderBuffer_2_valid ? _GEN_339 : _GEN_331; // @[LoadStoreQueue.scala 109:20]
  wire  _GEN_348 = io_reorderBuffer_2_valid ? _GEN_340 : _GEN_332; // @[LoadStoreQueue.scala 109:20]
  wire  _GEN_349 = io_reorderBuffer_2_valid ? _GEN_341 : _GEN_333; // @[LoadStoreQueue.scala 109:20]
  wire  _GEN_350 = io_reorderBuffer_2_valid ? _GEN_342 : _GEN_334; // @[LoadStoreQueue.scala 109:20]
  wire  _GEN_351 = io_reorderBuffer_2_valid ? _GEN_343 : _GEN_335; // @[LoadStoreQueue.scala 109:20]
  wire  _T_203 = io_reorderBuffer_3_bits_destinationTag_id == buffer_0_addressAndLoadResultTag_id &
    io_reorderBuffer_3_bits_destinationTag_threadId == buffer_0_addressAndLoadResultTag_threadId; // @[Tag.scala 13:25]
  wire  _T_204 = buffer_0_valid & _T_203; // @[LoadStoreQueue.scala 112:21]
  wire  _GEN_352 = _T_204 | _GEN_344; // @[LoadStoreQueue.scala 113:11 114:32]
  wire  _T_207 = io_reorderBuffer_3_bits_destinationTag_id == buffer_1_addressAndLoadResultTag_id &
    io_reorderBuffer_3_bits_destinationTag_threadId == buffer_1_addressAndLoadResultTag_threadId; // @[Tag.scala 13:25]
  wire  _T_208 = buffer_1_valid & _T_207; // @[LoadStoreQueue.scala 112:21]
  wire  _GEN_353 = _T_208 | _GEN_345; // @[LoadStoreQueue.scala 113:11 114:32]
  wire  _T_211 = io_reorderBuffer_3_bits_destinationTag_id == buffer_2_addressAndLoadResultTag_id &
    io_reorderBuffer_3_bits_destinationTag_threadId == buffer_2_addressAndLoadResultTag_threadId; // @[Tag.scala 13:25]
  wire  _T_212 = buffer_2_valid & _T_211; // @[LoadStoreQueue.scala 112:21]
  wire  _GEN_354 = _T_212 | _GEN_346; // @[LoadStoreQueue.scala 113:11 114:32]
  wire  _T_215 = io_reorderBuffer_3_bits_destinationTag_id == buffer_3_addressAndLoadResultTag_id &
    io_reorderBuffer_3_bits_destinationTag_threadId == buffer_3_addressAndLoadResultTag_threadId; // @[Tag.scala 13:25]
  wire  _T_216 = buffer_3_valid & _T_215; // @[LoadStoreQueue.scala 112:21]
  wire  _GEN_355 = _T_216 | _GEN_347; // @[LoadStoreQueue.scala 113:11 114:32]
  wire  _T_219 = io_reorderBuffer_3_bits_destinationTag_id == buffer_4_addressAndLoadResultTag_id &
    io_reorderBuffer_3_bits_destinationTag_threadId == buffer_4_addressAndLoadResultTag_threadId; // @[Tag.scala 13:25]
  wire  _T_220 = buffer_4_valid & _T_219; // @[LoadStoreQueue.scala 112:21]
  wire  _GEN_356 = _T_220 | _GEN_348; // @[LoadStoreQueue.scala 113:11 114:32]
  wire  _T_223 = io_reorderBuffer_3_bits_destinationTag_id == buffer_5_addressAndLoadResultTag_id &
    io_reorderBuffer_3_bits_destinationTag_threadId == buffer_5_addressAndLoadResultTag_threadId; // @[Tag.scala 13:25]
  wire  _T_224 = buffer_5_valid & _T_223; // @[LoadStoreQueue.scala 112:21]
  wire  _GEN_357 = _T_224 | _GEN_349; // @[LoadStoreQueue.scala 113:11 114:32]
  wire  _T_227 = io_reorderBuffer_3_bits_destinationTag_id == buffer_6_addressAndLoadResultTag_id &
    io_reorderBuffer_3_bits_destinationTag_threadId == buffer_6_addressAndLoadResultTag_threadId; // @[Tag.scala 13:25]
  wire  _T_228 = buffer_6_valid & _T_227; // @[LoadStoreQueue.scala 112:21]
  wire  _GEN_358 = _T_228 | _GEN_350; // @[LoadStoreQueue.scala 113:11 114:32]
  wire  _T_231 = io_reorderBuffer_3_bits_destinationTag_id == buffer_7_addressAndLoadResultTag_id &
    io_reorderBuffer_3_bits_destinationTag_threadId == buffer_7_addressAndLoadResultTag_threadId; // @[Tag.scala 13:25]
  wire  _T_232 = buffer_7_valid & _T_231; // @[LoadStoreQueue.scala 112:21]
  wire  _GEN_359 = _T_232 | _GEN_351; // @[LoadStoreQueue.scala 113:11 114:32]
  wire  _GEN_360 = io_reorderBuffer_3_valid ? _GEN_352 : _GEN_344; // @[LoadStoreQueue.scala 109:20]
  wire  _GEN_361 = io_reorderBuffer_3_valid ? _GEN_353 : _GEN_345; // @[LoadStoreQueue.scala 109:20]
  wire  _GEN_362 = io_reorderBuffer_3_valid ? _GEN_354 : _GEN_346; // @[LoadStoreQueue.scala 109:20]
  wire  _GEN_363 = io_reorderBuffer_3_valid ? _GEN_355 : _GEN_347; // @[LoadStoreQueue.scala 109:20]
  wire  _GEN_364 = io_reorderBuffer_3_valid ? _GEN_356 : _GEN_348; // @[LoadStoreQueue.scala 109:20]
  wire  _GEN_365 = io_reorderBuffer_3_valid ? _GEN_357 : _GEN_349; // @[LoadStoreQueue.scala 109:20]
  wire  _GEN_366 = io_reorderBuffer_3_valid ? _GEN_358 : _GEN_350; // @[LoadStoreQueue.scala 109:20]
  wire  _GEN_367 = io_reorderBuffer_3_valid ? _GEN_359 : _GEN_351; // @[LoadStoreQueue.scala 109:20]
  wire [3:0] _checkIndex_T = {{1'd0}, nextTail}; // @[LoadStoreQueue.scala 148:27]
  wire [2:0] checkIndex = _checkIndex_T[2:0]; // @[LoadStoreQueue.scala 148:27]
  wire  _GEN_369 = 3'h1 == checkIndex ? buffer_1_valid : buffer_0_valid; // @[LoadStoreQueue.scala 150:{36,36}]
  wire  _GEN_370 = 3'h2 == checkIndex ? buffer_2_valid : _GEN_369; // @[LoadStoreQueue.scala 150:{36,36}]
  wire  _GEN_371 = 3'h3 == checkIndex ? buffer_3_valid : _GEN_370; // @[LoadStoreQueue.scala 150:{36,36}]
  wire  _GEN_372 = 3'h4 == checkIndex ? buffer_4_valid : _GEN_371; // @[LoadStoreQueue.scala 150:{36,36}]
  wire  _GEN_373 = 3'h5 == checkIndex ? buffer_5_valid : _GEN_372; // @[LoadStoreQueue.scala 150:{36,36}]
  wire  _GEN_374 = 3'h6 == checkIndex ? buffer_6_valid : _GEN_373; // @[LoadStoreQueue.scala 150:{36,36}]
  wire  EntryValid_0 = 3'h7 == checkIndex ? buffer_7_valid : _GEN_374; // @[LoadStoreQueue.scala 150:{36,36}]
  wire [63:0] _GEN_377 = 3'h1 == checkIndex ? buffer_1_address : buffer_0_address; // @[LoadStoreQueue.scala 151:{18,18}]
  wire [63:0] _GEN_378 = 3'h2 == checkIndex ? buffer_2_address : _GEN_377; // @[LoadStoreQueue.scala 151:{18,18}]
  wire [63:0] _GEN_379 = 3'h3 == checkIndex ? buffer_3_address : _GEN_378; // @[LoadStoreQueue.scala 151:{18,18}]
  wire [63:0] _GEN_380 = 3'h4 == checkIndex ? buffer_4_address : _GEN_379; // @[LoadStoreQueue.scala 151:{18,18}]
  wire [63:0] _GEN_381 = 3'h5 == checkIndex ? buffer_5_address : _GEN_380; // @[LoadStoreQueue.scala 151:{18,18}]
  wire [63:0] _GEN_382 = 3'h6 == checkIndex ? buffer_6_address : _GEN_381; // @[LoadStoreQueue.scala 151:{18,18}]
  wire [63:0] _GEN_383 = 3'h7 == checkIndex ? buffer_7_address : _GEN_382; // @[LoadStoreQueue.scala 151:{18,18}]
  wire  _GEN_385 = 3'h1 == checkIndex ? buffer_1_addressValid : buffer_0_addressValid; // @[LoadStoreQueue.scala 152:{23,23}]
  wire  _GEN_386 = 3'h2 == checkIndex ? buffer_2_addressValid : _GEN_385; // @[LoadStoreQueue.scala 152:{23,23}]
  wire  _GEN_387 = 3'h3 == checkIndex ? buffer_3_addressValid : _GEN_386; // @[LoadStoreQueue.scala 152:{23,23}]
  wire  _GEN_388 = 3'h4 == checkIndex ? buffer_4_addressValid : _GEN_387; // @[LoadStoreQueue.scala 152:{23,23}]
  wire  _GEN_389 = 3'h5 == checkIndex ? buffer_5_addressValid : _GEN_388; // @[LoadStoreQueue.scala 152:{23,23}]
  wire  _GEN_390 = 3'h6 == checkIndex ? buffer_6_addressValid : _GEN_389; // @[LoadStoreQueue.scala 152:{23,23}]
  wire  _GEN_391 = 3'h7 == checkIndex ? buffer_7_addressValid : _GEN_390; // @[LoadStoreQueue.scala 152:{23,23}]
  wire  _checkOk_T = head != nextTail; // @[LoadStoreQueue.scala 171:24]
  wire  _checkOk_T_2 = head != nextTail & EntryValid_0 & _GEN_391; // @[LoadStoreQueue.scala 171:62]
  wire  _GEN_393 = 3'h1 == checkIndex ? buffer_1_info_accessType : buffer_0_info_accessType; // @[LoadStoreQueue.scala 174:{46,46}]
  wire  _GEN_394 = 3'h2 == checkIndex ? buffer_2_info_accessType : _GEN_393; // @[LoadStoreQueue.scala 174:{46,46}]
  wire  _GEN_395 = 3'h3 == checkIndex ? buffer_3_info_accessType : _GEN_394; // @[LoadStoreQueue.scala 174:{46,46}]
  wire  _GEN_396 = 3'h4 == checkIndex ? buffer_4_info_accessType : _GEN_395; // @[LoadStoreQueue.scala 174:{46,46}]
  wire  _GEN_397 = 3'h5 == checkIndex ? buffer_5_info_accessType : _GEN_396; // @[LoadStoreQueue.scala 174:{46,46}]
  wire  _GEN_398 = 3'h6 == checkIndex ? buffer_6_info_accessType : _GEN_397; // @[LoadStoreQueue.scala 174:{46,46}]
  wire  _GEN_399 = 3'h7 == checkIndex ? buffer_7_info_accessType : _GEN_398; // @[LoadStoreQueue.scala 174:{46,46}]
  wire  _GEN_401 = 3'h1 == checkIndex ? buffer_1_storeDataValid : buffer_0_storeDataValid; // @[LoadStoreQueue.scala 175:{57,57}]
  wire  _GEN_402 = 3'h2 == checkIndex ? buffer_2_storeDataValid : _GEN_401; // @[LoadStoreQueue.scala 175:{57,57}]
  wire  _GEN_403 = 3'h3 == checkIndex ? buffer_3_storeDataValid : _GEN_402; // @[LoadStoreQueue.scala 175:{57,57}]
  wire  _GEN_404 = 3'h4 == checkIndex ? buffer_4_storeDataValid : _GEN_403; // @[LoadStoreQueue.scala 175:{57,57}]
  wire  _GEN_405 = 3'h5 == checkIndex ? buffer_5_storeDataValid : _GEN_404; // @[LoadStoreQueue.scala 175:{57,57}]
  wire  _GEN_406 = 3'h6 == checkIndex ? buffer_6_storeDataValid : _GEN_405; // @[LoadStoreQueue.scala 175:{57,57}]
  wire  _GEN_407 = 3'h7 == checkIndex ? buffer_7_storeDataValid : _GEN_406; // @[LoadStoreQueue.scala 175:{57,57}]
  wire  _checkOk_T_7 = ~_GEN_399 & _GEN_407; // @[LoadStoreQueue.scala 175:57]
  wire  _GEN_409 = 3'h1 == checkIndex ? buffer_1_readyReorderSign : buffer_0_readyReorderSign; // @[LoadStoreQueue.scala 177:{28,28}]
  wire  _GEN_410 = 3'h2 == checkIndex ? buffer_2_readyReorderSign : _GEN_409; // @[LoadStoreQueue.scala 177:{28,28}]
  wire  _GEN_411 = 3'h3 == checkIndex ? buffer_3_readyReorderSign : _GEN_410; // @[LoadStoreQueue.scala 177:{28,28}]
  wire  _GEN_412 = 3'h4 == checkIndex ? buffer_4_readyReorderSign : _GEN_411; // @[LoadStoreQueue.scala 177:{28,28}]
  wire  _GEN_413 = 3'h5 == checkIndex ? buffer_5_readyReorderSign : _GEN_412; // @[LoadStoreQueue.scala 177:{28,28}]
  wire  _GEN_414 = 3'h6 == checkIndex ? buffer_6_readyReorderSign : _GEN_413; // @[LoadStoreQueue.scala 177:{28,28}]
  wire  _GEN_415 = 3'h7 == checkIndex ? buffer_7_readyReorderSign : _GEN_414; // @[LoadStoreQueue.scala 177:{28,28}]
  wire  _checkOk_T_8 = _checkOk_T_7 & _GEN_415; // @[LoadStoreQueue.scala 177:28]
  wire  _checkOk_T_9 = _GEN_399 | _checkOk_T_8; // @[LoadStoreQueue.scala 174:71]
  wire  _checkOk_T_10 = _checkOk_T_2 & _checkOk_T_9; // @[LoadStoreQueue.scala 173:22]
  wire  checkOk = EntryValid_0 & _checkOk_T_10; // @[LoadStoreQueue.scala 150:36 171:15 149:30]
  wire  _GEN_417 = 3'h1 == checkIndex ? buffer_1_addressAndLoadResultTag_threadId :
    buffer_0_addressAndLoadResultTag_threadId; // @[LoadStoreQueue.scala 182:{28,28}]
  wire  _GEN_418 = 3'h2 == checkIndex ? buffer_2_addressAndLoadResultTag_threadId : _GEN_417; // @[LoadStoreQueue.scala 182:{28,28}]
  wire  _GEN_419 = 3'h3 == checkIndex ? buffer_3_addressAndLoadResultTag_threadId : _GEN_418; // @[LoadStoreQueue.scala 182:{28,28}]
  wire  _GEN_420 = 3'h4 == checkIndex ? buffer_4_addressAndLoadResultTag_threadId : _GEN_419; // @[LoadStoreQueue.scala 182:{28,28}]
  wire  _GEN_421 = 3'h5 == checkIndex ? buffer_5_addressAndLoadResultTag_threadId : _GEN_420; // @[LoadStoreQueue.scala 182:{28,28}]
  wire  _GEN_422 = 3'h6 == checkIndex ? buffer_6_addressAndLoadResultTag_threadId : _GEN_421; // @[LoadStoreQueue.scala 182:{28,28}]
  wire  _GEN_423 = 3'h7 == checkIndex ? buffer_7_addressAndLoadResultTag_threadId : _GEN_422; // @[LoadStoreQueue.scala 182:{28,28}]
  wire [3:0] _GEN_425 = 3'h1 == checkIndex ? buffer_1_addressAndLoadResultTag_id : buffer_0_addressAndLoadResultTag_id; // @[LoadStoreQueue.scala 182:{28,28}]
  wire [3:0] _GEN_426 = 3'h2 == checkIndex ? buffer_2_addressAndLoadResultTag_id : _GEN_425; // @[LoadStoreQueue.scala 182:{28,28}]
  wire [3:0] _GEN_427 = 3'h3 == checkIndex ? buffer_3_addressAndLoadResultTag_id : _GEN_426; // @[LoadStoreQueue.scala 182:{28,28}]
  wire [3:0] _GEN_428 = 3'h4 == checkIndex ? buffer_4_addressAndLoadResultTag_id : _GEN_427; // @[LoadStoreQueue.scala 182:{28,28}]
  wire [3:0] _GEN_429 = 3'h5 == checkIndex ? buffer_5_addressAndLoadResultTag_id : _GEN_428; // @[LoadStoreQueue.scala 182:{28,28}]
  wire [3:0] _GEN_430 = 3'h6 == checkIndex ? buffer_6_addressAndLoadResultTag_id : _GEN_429; // @[LoadStoreQueue.scala 182:{28,28}]
  wire [3:0] _GEN_431 = 3'h7 == checkIndex ? buffer_7_addressAndLoadResultTag_id : _GEN_430; // @[LoadStoreQueue.scala 182:{28,28}]
  wire [63:0] _GEN_433 = 3'h1 == checkIndex ? buffer_1_storeData : buffer_0_storeData; // @[LoadStoreQueue.scala 183:{29,29}]
  wire [63:0] _GEN_434 = 3'h2 == checkIndex ? buffer_2_storeData : _GEN_433; // @[LoadStoreQueue.scala 183:{29,29}]
  wire [63:0] _GEN_435 = 3'h3 == checkIndex ? buffer_3_storeData : _GEN_434; // @[LoadStoreQueue.scala 183:{29,29}]
  wire [63:0] _GEN_436 = 3'h4 == checkIndex ? buffer_4_storeData : _GEN_435; // @[LoadStoreQueue.scala 183:{29,29}]
  wire [63:0] _GEN_437 = 3'h5 == checkIndex ? buffer_5_storeData : _GEN_436; // @[LoadStoreQueue.scala 183:{29,29}]
  wire [63:0] _GEN_438 = 3'h6 == checkIndex ? buffer_6_storeData : _GEN_437; // @[LoadStoreQueue.scala 183:{29,29}]
  wire [63:0] _GEN_439 = 3'h7 == checkIndex ? buffer_7_storeData : _GEN_438; // @[LoadStoreQueue.scala 183:{29,29}]
  wire  _GEN_441 = 3'h1 == checkIndex ? buffer_1_info_signed : buffer_0_info_signed; // @[LoadStoreQueue.scala 185:{35,35}]
  wire  _GEN_442 = 3'h2 == checkIndex ? buffer_2_info_signed : _GEN_441; // @[LoadStoreQueue.scala 185:{35,35}]
  wire  _GEN_443 = 3'h3 == checkIndex ? buffer_3_info_signed : _GEN_442; // @[LoadStoreQueue.scala 185:{35,35}]
  wire  _GEN_444 = 3'h4 == checkIndex ? buffer_4_info_signed : _GEN_443; // @[LoadStoreQueue.scala 185:{35,35}]
  wire  _GEN_445 = 3'h5 == checkIndex ? buffer_5_info_signed : _GEN_444; // @[LoadStoreQueue.scala 185:{35,35}]
  wire  _GEN_446 = 3'h6 == checkIndex ? buffer_6_info_signed : _GEN_445; // @[LoadStoreQueue.scala 185:{35,35}]
  wire  _GEN_447 = 3'h7 == checkIndex ? buffer_7_info_signed : _GEN_446; // @[LoadStoreQueue.scala 185:{35,35}]
  wire [1:0] _GEN_449 = 3'h1 == checkIndex ? buffer_1_info_accessWidth : buffer_0_info_accessWidth; // @[LoadStoreQueue.scala 185:{35,35}]
  wire [1:0] _GEN_450 = 3'h2 == checkIndex ? buffer_2_info_accessWidth : _GEN_449; // @[LoadStoreQueue.scala 185:{35,35}]
  wire [1:0] _GEN_451 = 3'h3 == checkIndex ? buffer_3_info_accessWidth : _GEN_450; // @[LoadStoreQueue.scala 185:{35,35}]
  wire [1:0] _GEN_452 = 3'h4 == checkIndex ? buffer_4_info_accessWidth : _GEN_451; // @[LoadStoreQueue.scala 185:{35,35}]
  wire [1:0] _GEN_453 = 3'h5 == checkIndex ? buffer_5_info_accessWidth : _GEN_452; // @[LoadStoreQueue.scala 185:{35,35}]
  wire [1:0] _GEN_454 = 3'h6 == checkIndex ? buffer_6_info_accessWidth : _GEN_453; // @[LoadStoreQueue.scala 185:{35,35}]
  wire [1:0] _GEN_455 = 3'h7 == checkIndex ? buffer_7_info_accessWidth : _GEN_454; // @[LoadStoreQueue.scala 185:{35,35}]
  wire  _GEN_456 = 3'h0 == checkIndex ? 1'h0 : _GEN_104; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_457 = 3'h1 == checkIndex ? 1'h0 : _GEN_105; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_458 = 3'h2 == checkIndex ? 1'h0 : _GEN_106; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_459 = 3'h3 == checkIndex ? 1'h0 : _GEN_107; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_460 = 3'h4 == checkIndex ? 1'h0 : _GEN_108; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_461 = 3'h5 == checkIndex ? 1'h0 : _GEN_109; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_462 = 3'h6 == checkIndex ? 1'h0 : _GEN_110; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_463 = 3'h7 == checkIndex ? 1'h0 : _GEN_111; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_464 = 3'h0 == checkIndex ? 1'h0 : _GEN_360; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_465 = 3'h1 == checkIndex ? 1'h0 : _GEN_361; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_466 = 3'h2 == checkIndex ? 1'h0 : _GEN_362; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_467 = 3'h3 == checkIndex ? 1'h0 : _GEN_363; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_468 = 3'h4 == checkIndex ? 1'h0 : _GEN_364; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_469 = 3'h5 == checkIndex ? 1'h0 : _GEN_365; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_470 = 3'h6 == checkIndex ? 1'h0 : _GEN_366; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_471 = 3'h7 == checkIndex ? 1'h0 : _GEN_367; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_472 = 3'h0 == checkIndex ? 1'h0 : _GEN_120; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_473 = 3'h1 == checkIndex ? 1'h0 : _GEN_121; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_474 = 3'h2 == checkIndex ? 1'h0 : _GEN_122; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_475 = 3'h3 == checkIndex ? 1'h0 : _GEN_123; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_476 = 3'h4 == checkIndex ? 1'h0 : _GEN_124; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_477 = 3'h5 == checkIndex ? 1'h0 : _GEN_125; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_478 = 3'h6 == checkIndex ? 1'h0 : _GEN_126; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_479 = 3'h7 == checkIndex ? 1'h0 : _GEN_127; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_480 = 3'h0 == checkIndex ? 1'h0 : _GEN_128; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_481 = 3'h1 == checkIndex ? 1'h0 : _GEN_129; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_482 = 3'h2 == checkIndex ? 1'h0 : _GEN_130; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_483 = 3'h3 == checkIndex ? 1'h0 : _GEN_131; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_484 = 3'h4 == checkIndex ? 1'h0 : _GEN_132; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_485 = 3'h5 == checkIndex ? 1'h0 : _GEN_133; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_486 = 3'h6 == checkIndex ? 1'h0 : _GEN_134; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_487 = 3'h7 == checkIndex ? 1'h0 : _GEN_135; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [1:0] _GEN_488 = 3'h0 == checkIndex ? 2'h0 : _GEN_136; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [1:0] _GEN_489 = 3'h1 == checkIndex ? 2'h0 : _GEN_137; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [1:0] _GEN_490 = 3'h2 == checkIndex ? 2'h0 : _GEN_138; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [1:0] _GEN_491 = 3'h3 == checkIndex ? 2'h0 : _GEN_139; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [1:0] _GEN_492 = 3'h4 == checkIndex ? 2'h0 : _GEN_140; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [1:0] _GEN_493 = 3'h5 == checkIndex ? 2'h0 : _GEN_141; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [1:0] _GEN_494 = 3'h6 == checkIndex ? 2'h0 : _GEN_142; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [1:0] _GEN_495 = 3'h7 == checkIndex ? 2'h0 : _GEN_143; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_496 = 3'h0 == checkIndex ? 1'h0 : _GEN_144; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_497 = 3'h1 == checkIndex ? 1'h0 : _GEN_145; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_498 = 3'h2 == checkIndex ? 1'h0 : _GEN_146; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_499 = 3'h3 == checkIndex ? 1'h0 : _GEN_147; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_500 = 3'h4 == checkIndex ? 1'h0 : _GEN_148; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_501 = 3'h5 == checkIndex ? 1'h0 : _GEN_149; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_502 = 3'h6 == checkIndex ? 1'h0 : _GEN_150; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_503 = 3'h7 == checkIndex ? 1'h0 : _GEN_151; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [3:0] _GEN_504 = 3'h0 == checkIndex ? 4'h0 : _GEN_152; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [3:0] _GEN_505 = 3'h1 == checkIndex ? 4'h0 : _GEN_153; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [3:0] _GEN_506 = 3'h2 == checkIndex ? 4'h0 : _GEN_154; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [3:0] _GEN_507 = 3'h3 == checkIndex ? 4'h0 : _GEN_155; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [3:0] _GEN_508 = 3'h4 == checkIndex ? 4'h0 : _GEN_156; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [3:0] _GEN_509 = 3'h5 == checkIndex ? 4'h0 : _GEN_157; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [3:0] _GEN_510 = 3'h6 == checkIndex ? 4'h0 : _GEN_158; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [3:0] _GEN_511 = 3'h7 == checkIndex ? 4'h0 : _GEN_159; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [63:0] _GEN_512 = 3'h0 == checkIndex ? 64'h0 : _GEN_216; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [63:0] _GEN_513 = 3'h1 == checkIndex ? 64'h0 : _GEN_228; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [63:0] _GEN_514 = 3'h2 == checkIndex ? 64'h0 : _GEN_240; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [63:0] _GEN_515 = 3'h3 == checkIndex ? 64'h0 : _GEN_252; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [63:0] _GEN_516 = 3'h4 == checkIndex ? 64'h0 : _GEN_264; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [63:0] _GEN_517 = 3'h5 == checkIndex ? 64'h0 : _GEN_276; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [63:0] _GEN_518 = 3'h6 == checkIndex ? 64'h0 : _GEN_288; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [63:0] _GEN_519 = 3'h7 == checkIndex ? 64'h0 : _GEN_300; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_520 = 3'h0 == checkIndex ? 1'h0 : _GEN_217; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_521 = 3'h1 == checkIndex ? 1'h0 : _GEN_229; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_522 = 3'h2 == checkIndex ? 1'h0 : _GEN_241; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_523 = 3'h3 == checkIndex ? 1'h0 : _GEN_253; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_524 = 3'h4 == checkIndex ? 1'h0 : _GEN_265; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_525 = 3'h5 == checkIndex ? 1'h0 : _GEN_277; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_526 = 3'h6 == checkIndex ? 1'h0 : _GEN_289; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_527 = 3'h7 == checkIndex ? 1'h0 : _GEN_301; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_528 = 3'h0 == checkIndex ? 1'h0 : _GEN_176; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_529 = 3'h1 == checkIndex ? 1'h0 : _GEN_177; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_530 = 3'h2 == checkIndex ? 1'h0 : _GEN_178; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_531 = 3'h3 == checkIndex ? 1'h0 : _GEN_179; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_532 = 3'h4 == checkIndex ? 1'h0 : _GEN_180; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_533 = 3'h5 == checkIndex ? 1'h0 : _GEN_181; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_534 = 3'h6 == checkIndex ? 1'h0 : _GEN_182; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_535 = 3'h7 == checkIndex ? 1'h0 : _GEN_183; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [3:0] _GEN_536 = 3'h0 == checkIndex ? 4'h0 : _GEN_184; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [3:0] _GEN_537 = 3'h1 == checkIndex ? 4'h0 : _GEN_185; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [3:0] _GEN_538 = 3'h2 == checkIndex ? 4'h0 : _GEN_186; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [3:0] _GEN_539 = 3'h3 == checkIndex ? 4'h0 : _GEN_187; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [3:0] _GEN_540 = 3'h4 == checkIndex ? 4'h0 : _GEN_188; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [3:0] _GEN_541 = 3'h5 == checkIndex ? 4'h0 : _GEN_189; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [3:0] _GEN_542 = 3'h6 == checkIndex ? 4'h0 : _GEN_190; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [3:0] _GEN_543 = 3'h7 == checkIndex ? 4'h0 : _GEN_191; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [63:0] _GEN_544 = 3'h0 == checkIndex ? 64'h0 : _GEN_218; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [63:0] _GEN_545 = 3'h1 == checkIndex ? 64'h0 : _GEN_230; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [63:0] _GEN_546 = 3'h2 == checkIndex ? 64'h0 : _GEN_242; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [63:0] _GEN_547 = 3'h3 == checkIndex ? 64'h0 : _GEN_254; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [63:0] _GEN_548 = 3'h4 == checkIndex ? 64'h0 : _GEN_266; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [63:0] _GEN_549 = 3'h5 == checkIndex ? 64'h0 : _GEN_278; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [63:0] _GEN_550 = 3'h6 == checkIndex ? 64'h0 : _GEN_290; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [63:0] _GEN_551 = 3'h7 == checkIndex ? 64'h0 : _GEN_302; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_552 = 3'h0 == checkIndex ? 1'h0 : _GEN_219; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_553 = 3'h1 == checkIndex ? 1'h0 : _GEN_231; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_554 = 3'h2 == checkIndex ? 1'h0 : _GEN_243; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_555 = 3'h3 == checkIndex ? 1'h0 : _GEN_255; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_556 = 3'h4 == checkIndex ? 1'h0 : _GEN_267; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_557 = 3'h5 == checkIndex ? 1'h0 : _GEN_279; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_558 = 3'h6 == checkIndex ? 1'h0 : _GEN_291; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_559 = 3'h7 == checkIndex ? 1'h0 : _GEN_303; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_560 = io_memory_ready ? _GEN_456 : _GEN_104; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_561 = io_memory_ready ? _GEN_457 : _GEN_105; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_562 = io_memory_ready ? _GEN_458 : _GEN_106; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_563 = io_memory_ready ? _GEN_459 : _GEN_107; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_564 = io_memory_ready ? _GEN_460 : _GEN_108; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_565 = io_memory_ready ? _GEN_461 : _GEN_109; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_566 = io_memory_ready ? _GEN_462 : _GEN_110; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_567 = io_memory_ready ? _GEN_463 : _GEN_111; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_568 = io_memory_ready ? _GEN_464 : _GEN_360; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_569 = io_memory_ready ? _GEN_465 : _GEN_361; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_570 = io_memory_ready ? _GEN_466 : _GEN_362; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_571 = io_memory_ready ? _GEN_467 : _GEN_363; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_572 = io_memory_ready ? _GEN_468 : _GEN_364; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_573 = io_memory_ready ? _GEN_469 : _GEN_365; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_574 = io_memory_ready ? _GEN_470 : _GEN_366; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_575 = io_memory_ready ? _GEN_471 : _GEN_367; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_576 = io_memory_ready ? _GEN_472 : _GEN_120; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_577 = io_memory_ready ? _GEN_473 : _GEN_121; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_578 = io_memory_ready ? _GEN_474 : _GEN_122; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_579 = io_memory_ready ? _GEN_475 : _GEN_123; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_580 = io_memory_ready ? _GEN_476 : _GEN_124; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_581 = io_memory_ready ? _GEN_477 : _GEN_125; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_582 = io_memory_ready ? _GEN_478 : _GEN_126; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_583 = io_memory_ready ? _GEN_479 : _GEN_127; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_584 = io_memory_ready ? _GEN_480 : _GEN_128; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_585 = io_memory_ready ? _GEN_481 : _GEN_129; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_586 = io_memory_ready ? _GEN_482 : _GEN_130; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_587 = io_memory_ready ? _GEN_483 : _GEN_131; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_588 = io_memory_ready ? _GEN_484 : _GEN_132; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_589 = io_memory_ready ? _GEN_485 : _GEN_133; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_590 = io_memory_ready ? _GEN_486 : _GEN_134; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_591 = io_memory_ready ? _GEN_487 : _GEN_135; // @[LoadStoreQueue.scala 186:31]
  wire [1:0] _GEN_592 = io_memory_ready ? _GEN_488 : _GEN_136; // @[LoadStoreQueue.scala 186:31]
  wire [1:0] _GEN_593 = io_memory_ready ? _GEN_489 : _GEN_137; // @[LoadStoreQueue.scala 186:31]
  wire [1:0] _GEN_594 = io_memory_ready ? _GEN_490 : _GEN_138; // @[LoadStoreQueue.scala 186:31]
  wire [1:0] _GEN_595 = io_memory_ready ? _GEN_491 : _GEN_139; // @[LoadStoreQueue.scala 186:31]
  wire [1:0] _GEN_596 = io_memory_ready ? _GEN_492 : _GEN_140; // @[LoadStoreQueue.scala 186:31]
  wire [1:0] _GEN_597 = io_memory_ready ? _GEN_493 : _GEN_141; // @[LoadStoreQueue.scala 186:31]
  wire [1:0] _GEN_598 = io_memory_ready ? _GEN_494 : _GEN_142; // @[LoadStoreQueue.scala 186:31]
  wire [1:0] _GEN_599 = io_memory_ready ? _GEN_495 : _GEN_143; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_600 = io_memory_ready ? _GEN_496 : _GEN_144; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_601 = io_memory_ready ? _GEN_497 : _GEN_145; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_602 = io_memory_ready ? _GEN_498 : _GEN_146; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_603 = io_memory_ready ? _GEN_499 : _GEN_147; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_604 = io_memory_ready ? _GEN_500 : _GEN_148; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_605 = io_memory_ready ? _GEN_501 : _GEN_149; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_606 = io_memory_ready ? _GEN_502 : _GEN_150; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_607 = io_memory_ready ? _GEN_503 : _GEN_151; // @[LoadStoreQueue.scala 186:31]
  wire [3:0] _GEN_608 = io_memory_ready ? _GEN_504 : _GEN_152; // @[LoadStoreQueue.scala 186:31]
  wire [3:0] _GEN_609 = io_memory_ready ? _GEN_505 : _GEN_153; // @[LoadStoreQueue.scala 186:31]
  wire [3:0] _GEN_610 = io_memory_ready ? _GEN_506 : _GEN_154; // @[LoadStoreQueue.scala 186:31]
  wire [3:0] _GEN_611 = io_memory_ready ? _GEN_507 : _GEN_155; // @[LoadStoreQueue.scala 186:31]
  wire [3:0] _GEN_612 = io_memory_ready ? _GEN_508 : _GEN_156; // @[LoadStoreQueue.scala 186:31]
  wire [3:0] _GEN_613 = io_memory_ready ? _GEN_509 : _GEN_157; // @[LoadStoreQueue.scala 186:31]
  wire [3:0] _GEN_614 = io_memory_ready ? _GEN_510 : _GEN_158; // @[LoadStoreQueue.scala 186:31]
  wire [3:0] _GEN_615 = io_memory_ready ? _GEN_511 : _GEN_159; // @[LoadStoreQueue.scala 186:31]
  wire [63:0] _GEN_616 = io_memory_ready ? _GEN_512 : _GEN_216; // @[LoadStoreQueue.scala 186:31]
  wire [63:0] _GEN_617 = io_memory_ready ? _GEN_513 : _GEN_228; // @[LoadStoreQueue.scala 186:31]
  wire [63:0] _GEN_618 = io_memory_ready ? _GEN_514 : _GEN_240; // @[LoadStoreQueue.scala 186:31]
  wire [63:0] _GEN_619 = io_memory_ready ? _GEN_515 : _GEN_252; // @[LoadStoreQueue.scala 186:31]
  wire [63:0] _GEN_620 = io_memory_ready ? _GEN_516 : _GEN_264; // @[LoadStoreQueue.scala 186:31]
  wire [63:0] _GEN_621 = io_memory_ready ? _GEN_517 : _GEN_276; // @[LoadStoreQueue.scala 186:31]
  wire [63:0] _GEN_622 = io_memory_ready ? _GEN_518 : _GEN_288; // @[LoadStoreQueue.scala 186:31]
  wire [63:0] _GEN_623 = io_memory_ready ? _GEN_519 : _GEN_300; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_624 = io_memory_ready ? _GEN_520 : _GEN_217; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_625 = io_memory_ready ? _GEN_521 : _GEN_229; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_626 = io_memory_ready ? _GEN_522 : _GEN_241; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_627 = io_memory_ready ? _GEN_523 : _GEN_253; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_628 = io_memory_ready ? _GEN_524 : _GEN_265; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_629 = io_memory_ready ? _GEN_525 : _GEN_277; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_630 = io_memory_ready ? _GEN_526 : _GEN_289; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_631 = io_memory_ready ? _GEN_527 : _GEN_301; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_632 = io_memory_ready ? _GEN_528 : _GEN_176; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_633 = io_memory_ready ? _GEN_529 : _GEN_177; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_634 = io_memory_ready ? _GEN_530 : _GEN_178; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_635 = io_memory_ready ? _GEN_531 : _GEN_179; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_636 = io_memory_ready ? _GEN_532 : _GEN_180; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_637 = io_memory_ready ? _GEN_533 : _GEN_181; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_638 = io_memory_ready ? _GEN_534 : _GEN_182; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_639 = io_memory_ready ? _GEN_535 : _GEN_183; // @[LoadStoreQueue.scala 186:31]
  wire [3:0] _GEN_640 = io_memory_ready ? _GEN_536 : _GEN_184; // @[LoadStoreQueue.scala 186:31]
  wire [3:0] _GEN_641 = io_memory_ready ? _GEN_537 : _GEN_185; // @[LoadStoreQueue.scala 186:31]
  wire [3:0] _GEN_642 = io_memory_ready ? _GEN_538 : _GEN_186; // @[LoadStoreQueue.scala 186:31]
  wire [3:0] _GEN_643 = io_memory_ready ? _GEN_539 : _GEN_187; // @[LoadStoreQueue.scala 186:31]
  wire [3:0] _GEN_644 = io_memory_ready ? _GEN_540 : _GEN_188; // @[LoadStoreQueue.scala 186:31]
  wire [3:0] _GEN_645 = io_memory_ready ? _GEN_541 : _GEN_189; // @[LoadStoreQueue.scala 186:31]
  wire [3:0] _GEN_646 = io_memory_ready ? _GEN_542 : _GEN_190; // @[LoadStoreQueue.scala 186:31]
  wire [3:0] _GEN_647 = io_memory_ready ? _GEN_543 : _GEN_191; // @[LoadStoreQueue.scala 186:31]
  wire [63:0] _GEN_648 = io_memory_ready ? _GEN_544 : _GEN_218; // @[LoadStoreQueue.scala 186:31]
  wire [63:0] _GEN_649 = io_memory_ready ? _GEN_545 : _GEN_230; // @[LoadStoreQueue.scala 186:31]
  wire [63:0] _GEN_650 = io_memory_ready ? _GEN_546 : _GEN_242; // @[LoadStoreQueue.scala 186:31]
  wire [63:0] _GEN_651 = io_memory_ready ? _GEN_547 : _GEN_254; // @[LoadStoreQueue.scala 186:31]
  wire [63:0] _GEN_652 = io_memory_ready ? _GEN_548 : _GEN_266; // @[LoadStoreQueue.scala 186:31]
  wire [63:0] _GEN_653 = io_memory_ready ? _GEN_549 : _GEN_278; // @[LoadStoreQueue.scala 186:31]
  wire [63:0] _GEN_654 = io_memory_ready ? _GEN_550 : _GEN_290; // @[LoadStoreQueue.scala 186:31]
  wire [63:0] _GEN_655 = io_memory_ready ? _GEN_551 : _GEN_302; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_656 = io_memory_ready ? _GEN_552 : _GEN_219; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_657 = io_memory_ready ? _GEN_553 : _GEN_231; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_658 = io_memory_ready ? _GEN_554 : _GEN_243; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_659 = io_memory_ready ? _GEN_555 : _GEN_255; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_660 = io_memory_ready ? _GEN_556 : _GEN_267; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_661 = io_memory_ready ? _GEN_557 : _GEN_279; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_662 = io_memory_ready ? _GEN_558 : _GEN_291; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_663 = io_memory_ready ? _GEN_559 : _GEN_303; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_671 = checkOk ? _GEN_560 : _GEN_104; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_672 = checkOk ? _GEN_561 : _GEN_105; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_673 = checkOk ? _GEN_562 : _GEN_106; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_674 = checkOk ? _GEN_563 : _GEN_107; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_675 = checkOk ? _GEN_564 : _GEN_108; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_676 = checkOk ? _GEN_565 : _GEN_109; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_677 = checkOk ? _GEN_566 : _GEN_110; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_678 = checkOk ? _GEN_567 : _GEN_111; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_679 = checkOk ? _GEN_568 : _GEN_360; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_680 = checkOk ? _GEN_569 : _GEN_361; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_681 = checkOk ? _GEN_570 : _GEN_362; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_682 = checkOk ? _GEN_571 : _GEN_363; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_683 = checkOk ? _GEN_572 : _GEN_364; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_684 = checkOk ? _GEN_573 : _GEN_365; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_685 = checkOk ? _GEN_574 : _GEN_366; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_686 = checkOk ? _GEN_575 : _GEN_367; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_687 = checkOk ? _GEN_576 : _GEN_120; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_688 = checkOk ? _GEN_577 : _GEN_121; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_689 = checkOk ? _GEN_578 : _GEN_122; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_690 = checkOk ? _GEN_579 : _GEN_123; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_691 = checkOk ? _GEN_580 : _GEN_124; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_692 = checkOk ? _GEN_581 : _GEN_125; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_693 = checkOk ? _GEN_582 : _GEN_126; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_694 = checkOk ? _GEN_583 : _GEN_127; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_695 = checkOk ? _GEN_584 : _GEN_128; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_696 = checkOk ? _GEN_585 : _GEN_129; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_697 = checkOk ? _GEN_586 : _GEN_130; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_698 = checkOk ? _GEN_587 : _GEN_131; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_699 = checkOk ? _GEN_588 : _GEN_132; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_700 = checkOk ? _GEN_589 : _GEN_133; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_701 = checkOk ? _GEN_590 : _GEN_134; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_702 = checkOk ? _GEN_591 : _GEN_135; // @[LoadStoreQueue.scala 181:31]
  wire [1:0] _GEN_703 = checkOk ? _GEN_592 : _GEN_136; // @[LoadStoreQueue.scala 181:31]
  wire [1:0] _GEN_704 = checkOk ? _GEN_593 : _GEN_137; // @[LoadStoreQueue.scala 181:31]
  wire [1:0] _GEN_705 = checkOk ? _GEN_594 : _GEN_138; // @[LoadStoreQueue.scala 181:31]
  wire [1:0] _GEN_706 = checkOk ? _GEN_595 : _GEN_139; // @[LoadStoreQueue.scala 181:31]
  wire [1:0] _GEN_707 = checkOk ? _GEN_596 : _GEN_140; // @[LoadStoreQueue.scala 181:31]
  wire [1:0] _GEN_708 = checkOk ? _GEN_597 : _GEN_141; // @[LoadStoreQueue.scala 181:31]
  wire [1:0] _GEN_709 = checkOk ? _GEN_598 : _GEN_142; // @[LoadStoreQueue.scala 181:31]
  wire [1:0] _GEN_710 = checkOk ? _GEN_599 : _GEN_143; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_711 = checkOk ? _GEN_600 : _GEN_144; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_712 = checkOk ? _GEN_601 : _GEN_145; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_713 = checkOk ? _GEN_602 : _GEN_146; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_714 = checkOk ? _GEN_603 : _GEN_147; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_715 = checkOk ? _GEN_604 : _GEN_148; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_716 = checkOk ? _GEN_605 : _GEN_149; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_717 = checkOk ? _GEN_606 : _GEN_150; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_718 = checkOk ? _GEN_607 : _GEN_151; // @[LoadStoreQueue.scala 181:31]
  wire [3:0] _GEN_719 = checkOk ? _GEN_608 : _GEN_152; // @[LoadStoreQueue.scala 181:31]
  wire [3:0] _GEN_720 = checkOk ? _GEN_609 : _GEN_153; // @[LoadStoreQueue.scala 181:31]
  wire [3:0] _GEN_721 = checkOk ? _GEN_610 : _GEN_154; // @[LoadStoreQueue.scala 181:31]
  wire [3:0] _GEN_722 = checkOk ? _GEN_611 : _GEN_155; // @[LoadStoreQueue.scala 181:31]
  wire [3:0] _GEN_723 = checkOk ? _GEN_612 : _GEN_156; // @[LoadStoreQueue.scala 181:31]
  wire [3:0] _GEN_724 = checkOk ? _GEN_613 : _GEN_157; // @[LoadStoreQueue.scala 181:31]
  wire [3:0] _GEN_725 = checkOk ? _GEN_614 : _GEN_158; // @[LoadStoreQueue.scala 181:31]
  wire [3:0] _GEN_726 = checkOk ? _GEN_615 : _GEN_159; // @[LoadStoreQueue.scala 181:31]
  wire [63:0] _GEN_727 = checkOk ? _GEN_616 : _GEN_216; // @[LoadStoreQueue.scala 181:31]
  wire [63:0] _GEN_728 = checkOk ? _GEN_617 : _GEN_228; // @[LoadStoreQueue.scala 181:31]
  wire [63:0] _GEN_729 = checkOk ? _GEN_618 : _GEN_240; // @[LoadStoreQueue.scala 181:31]
  wire [63:0] _GEN_730 = checkOk ? _GEN_619 : _GEN_252; // @[LoadStoreQueue.scala 181:31]
  wire [63:0] _GEN_731 = checkOk ? _GEN_620 : _GEN_264; // @[LoadStoreQueue.scala 181:31]
  wire [63:0] _GEN_732 = checkOk ? _GEN_621 : _GEN_276; // @[LoadStoreQueue.scala 181:31]
  wire [63:0] _GEN_733 = checkOk ? _GEN_622 : _GEN_288; // @[LoadStoreQueue.scala 181:31]
  wire [63:0] _GEN_734 = checkOk ? _GEN_623 : _GEN_300; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_735 = checkOk ? _GEN_624 : _GEN_217; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_736 = checkOk ? _GEN_625 : _GEN_229; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_737 = checkOk ? _GEN_626 : _GEN_241; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_738 = checkOk ? _GEN_627 : _GEN_253; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_739 = checkOk ? _GEN_628 : _GEN_265; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_740 = checkOk ? _GEN_629 : _GEN_277; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_741 = checkOk ? _GEN_630 : _GEN_289; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_742 = checkOk ? _GEN_631 : _GEN_301; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_743 = checkOk ? _GEN_632 : _GEN_176; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_744 = checkOk ? _GEN_633 : _GEN_177; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_745 = checkOk ? _GEN_634 : _GEN_178; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_746 = checkOk ? _GEN_635 : _GEN_179; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_747 = checkOk ? _GEN_636 : _GEN_180; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_748 = checkOk ? _GEN_637 : _GEN_181; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_749 = checkOk ? _GEN_638 : _GEN_182; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_750 = checkOk ? _GEN_639 : _GEN_183; // @[LoadStoreQueue.scala 181:31]
  wire [3:0] _GEN_751 = checkOk ? _GEN_640 : _GEN_184; // @[LoadStoreQueue.scala 181:31]
  wire [3:0] _GEN_752 = checkOk ? _GEN_641 : _GEN_185; // @[LoadStoreQueue.scala 181:31]
  wire [3:0] _GEN_753 = checkOk ? _GEN_642 : _GEN_186; // @[LoadStoreQueue.scala 181:31]
  wire [3:0] _GEN_754 = checkOk ? _GEN_643 : _GEN_187; // @[LoadStoreQueue.scala 181:31]
  wire [3:0] _GEN_755 = checkOk ? _GEN_644 : _GEN_188; // @[LoadStoreQueue.scala 181:31]
  wire [3:0] _GEN_756 = checkOk ? _GEN_645 : _GEN_189; // @[LoadStoreQueue.scala 181:31]
  wire [3:0] _GEN_757 = checkOk ? _GEN_646 : _GEN_190; // @[LoadStoreQueue.scala 181:31]
  wire [3:0] _GEN_758 = checkOk ? _GEN_647 : _GEN_191; // @[LoadStoreQueue.scala 181:31]
  wire [63:0] _GEN_759 = checkOk ? _GEN_648 : _GEN_218; // @[LoadStoreQueue.scala 181:31]
  wire [63:0] _GEN_760 = checkOk ? _GEN_649 : _GEN_230; // @[LoadStoreQueue.scala 181:31]
  wire [63:0] _GEN_761 = checkOk ? _GEN_650 : _GEN_242; // @[LoadStoreQueue.scala 181:31]
  wire [63:0] _GEN_762 = checkOk ? _GEN_651 : _GEN_254; // @[LoadStoreQueue.scala 181:31]
  wire [63:0] _GEN_763 = checkOk ? _GEN_652 : _GEN_266; // @[LoadStoreQueue.scala 181:31]
  wire [63:0] _GEN_764 = checkOk ? _GEN_653 : _GEN_278; // @[LoadStoreQueue.scala 181:31]
  wire [63:0] _GEN_765 = checkOk ? _GEN_654 : _GEN_290; // @[LoadStoreQueue.scala 181:31]
  wire [63:0] _GEN_766 = checkOk ? _GEN_655 : _GEN_302; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_767 = checkOk ? _GEN_656 : _GEN_219; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_768 = checkOk ? _GEN_657 : _GEN_231; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_769 = checkOk ? _GEN_658 : _GEN_243; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_770 = checkOk ? _GEN_659 : _GEN_255; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_771 = checkOk ? _GEN_660 : _GEN_267; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_772 = checkOk ? _GEN_661 : _GEN_279; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_773 = checkOk ? _GEN_662 : _GEN_291; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_774 = checkOk ? _GEN_663 : _GEN_303; // @[LoadStoreQueue.scala 181:31]
  wire [63:0] Address_0 = EntryValid_0 ? _GEN_383 : 64'h0; // @[LoadStoreQueue.scala 150:36 151:18 130:25]
  wire  AddressValid_0 = EntryValid_0 & _GEN_391; // @[LoadStoreQueue.scala 150:36 152:23 133:30]
  wire  _GEN_779 = EntryValid_0 & checkOk; // @[LoadStoreQueue.scala 146:19 150:36 179:23]
  wire  _GEN_787 = EntryValid_0 ? _GEN_671 : _GEN_104; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_788 = EntryValid_0 ? _GEN_672 : _GEN_105; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_789 = EntryValid_0 ? _GEN_673 : _GEN_106; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_790 = EntryValid_0 ? _GEN_674 : _GEN_107; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_791 = EntryValid_0 ? _GEN_675 : _GEN_108; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_792 = EntryValid_0 ? _GEN_676 : _GEN_109; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_793 = EntryValid_0 ? _GEN_677 : _GEN_110; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_794 = EntryValid_0 ? _GEN_678 : _GEN_111; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_795 = EntryValid_0 ? _GEN_679 : _GEN_360; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_796 = EntryValid_0 ? _GEN_680 : _GEN_361; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_797 = EntryValid_0 ? _GEN_681 : _GEN_362; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_798 = EntryValid_0 ? _GEN_682 : _GEN_363; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_799 = EntryValid_0 ? _GEN_683 : _GEN_364; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_800 = EntryValid_0 ? _GEN_684 : _GEN_365; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_801 = EntryValid_0 ? _GEN_685 : _GEN_366; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_802 = EntryValid_0 ? _GEN_686 : _GEN_367; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_803 = EntryValid_0 ? _GEN_687 : _GEN_120; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_804 = EntryValid_0 ? _GEN_688 : _GEN_121; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_805 = EntryValid_0 ? _GEN_689 : _GEN_122; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_806 = EntryValid_0 ? _GEN_690 : _GEN_123; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_807 = EntryValid_0 ? _GEN_691 : _GEN_124; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_808 = EntryValid_0 ? _GEN_692 : _GEN_125; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_809 = EntryValid_0 ? _GEN_693 : _GEN_126; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_810 = EntryValid_0 ? _GEN_694 : _GEN_127; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_811 = EntryValid_0 ? _GEN_695 : _GEN_128; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_812 = EntryValid_0 ? _GEN_696 : _GEN_129; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_813 = EntryValid_0 ? _GEN_697 : _GEN_130; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_814 = EntryValid_0 ? _GEN_698 : _GEN_131; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_815 = EntryValid_0 ? _GEN_699 : _GEN_132; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_816 = EntryValid_0 ? _GEN_700 : _GEN_133; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_817 = EntryValid_0 ? _GEN_701 : _GEN_134; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_818 = EntryValid_0 ? _GEN_702 : _GEN_135; // @[LoadStoreQueue.scala 150:36]
  wire [1:0] _GEN_819 = EntryValid_0 ? _GEN_703 : _GEN_136; // @[LoadStoreQueue.scala 150:36]
  wire [1:0] _GEN_820 = EntryValid_0 ? _GEN_704 : _GEN_137; // @[LoadStoreQueue.scala 150:36]
  wire [1:0] _GEN_821 = EntryValid_0 ? _GEN_705 : _GEN_138; // @[LoadStoreQueue.scala 150:36]
  wire [1:0] _GEN_822 = EntryValid_0 ? _GEN_706 : _GEN_139; // @[LoadStoreQueue.scala 150:36]
  wire [1:0] _GEN_823 = EntryValid_0 ? _GEN_707 : _GEN_140; // @[LoadStoreQueue.scala 150:36]
  wire [1:0] _GEN_824 = EntryValid_0 ? _GEN_708 : _GEN_141; // @[LoadStoreQueue.scala 150:36]
  wire [1:0] _GEN_825 = EntryValid_0 ? _GEN_709 : _GEN_142; // @[LoadStoreQueue.scala 150:36]
  wire [1:0] _GEN_826 = EntryValid_0 ? _GEN_710 : _GEN_143; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_827 = EntryValid_0 ? _GEN_711 : _GEN_144; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_828 = EntryValid_0 ? _GEN_712 : _GEN_145; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_829 = EntryValid_0 ? _GEN_713 : _GEN_146; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_830 = EntryValid_0 ? _GEN_714 : _GEN_147; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_831 = EntryValid_0 ? _GEN_715 : _GEN_148; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_832 = EntryValid_0 ? _GEN_716 : _GEN_149; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_833 = EntryValid_0 ? _GEN_717 : _GEN_150; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_834 = EntryValid_0 ? _GEN_718 : _GEN_151; // @[LoadStoreQueue.scala 150:36]
  wire [3:0] _GEN_835 = EntryValid_0 ? _GEN_719 : _GEN_152; // @[LoadStoreQueue.scala 150:36]
  wire [3:0] _GEN_836 = EntryValid_0 ? _GEN_720 : _GEN_153; // @[LoadStoreQueue.scala 150:36]
  wire [3:0] _GEN_837 = EntryValid_0 ? _GEN_721 : _GEN_154; // @[LoadStoreQueue.scala 150:36]
  wire [3:0] _GEN_838 = EntryValid_0 ? _GEN_722 : _GEN_155; // @[LoadStoreQueue.scala 150:36]
  wire [3:0] _GEN_839 = EntryValid_0 ? _GEN_723 : _GEN_156; // @[LoadStoreQueue.scala 150:36]
  wire [3:0] _GEN_840 = EntryValid_0 ? _GEN_724 : _GEN_157; // @[LoadStoreQueue.scala 150:36]
  wire [3:0] _GEN_841 = EntryValid_0 ? _GEN_725 : _GEN_158; // @[LoadStoreQueue.scala 150:36]
  wire [3:0] _GEN_842 = EntryValid_0 ? _GEN_726 : _GEN_159; // @[LoadStoreQueue.scala 150:36]
  wire [63:0] _GEN_843 = EntryValid_0 ? _GEN_727 : _GEN_216; // @[LoadStoreQueue.scala 150:36]
  wire [63:0] _GEN_844 = EntryValid_0 ? _GEN_728 : _GEN_228; // @[LoadStoreQueue.scala 150:36]
  wire [63:0] _GEN_845 = EntryValid_0 ? _GEN_729 : _GEN_240; // @[LoadStoreQueue.scala 150:36]
  wire [63:0] _GEN_846 = EntryValid_0 ? _GEN_730 : _GEN_252; // @[LoadStoreQueue.scala 150:36]
  wire [63:0] _GEN_847 = EntryValid_0 ? _GEN_731 : _GEN_264; // @[LoadStoreQueue.scala 150:36]
  wire [63:0] _GEN_848 = EntryValid_0 ? _GEN_732 : _GEN_276; // @[LoadStoreQueue.scala 150:36]
  wire [63:0] _GEN_849 = EntryValid_0 ? _GEN_733 : _GEN_288; // @[LoadStoreQueue.scala 150:36]
  wire [63:0] _GEN_850 = EntryValid_0 ? _GEN_734 : _GEN_300; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_851 = EntryValid_0 ? _GEN_735 : _GEN_217; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_852 = EntryValid_0 ? _GEN_736 : _GEN_229; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_853 = EntryValid_0 ? _GEN_737 : _GEN_241; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_854 = EntryValid_0 ? _GEN_738 : _GEN_253; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_855 = EntryValid_0 ? _GEN_739 : _GEN_265; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_856 = EntryValid_0 ? _GEN_740 : _GEN_277; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_857 = EntryValid_0 ? _GEN_741 : _GEN_289; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_858 = EntryValid_0 ? _GEN_742 : _GEN_301; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_859 = EntryValid_0 ? _GEN_743 : _GEN_176; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_860 = EntryValid_0 ? _GEN_744 : _GEN_177; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_861 = EntryValid_0 ? _GEN_745 : _GEN_178; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_862 = EntryValid_0 ? _GEN_746 : _GEN_179; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_863 = EntryValid_0 ? _GEN_747 : _GEN_180; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_864 = EntryValid_0 ? _GEN_748 : _GEN_181; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_865 = EntryValid_0 ? _GEN_749 : _GEN_182; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_866 = EntryValid_0 ? _GEN_750 : _GEN_183; // @[LoadStoreQueue.scala 150:36]
  wire [3:0] _GEN_867 = EntryValid_0 ? _GEN_751 : _GEN_184; // @[LoadStoreQueue.scala 150:36]
  wire [3:0] _GEN_868 = EntryValid_0 ? _GEN_752 : _GEN_185; // @[LoadStoreQueue.scala 150:36]
  wire [3:0] _GEN_869 = EntryValid_0 ? _GEN_753 : _GEN_186; // @[LoadStoreQueue.scala 150:36]
  wire [3:0] _GEN_870 = EntryValid_0 ? _GEN_754 : _GEN_187; // @[LoadStoreQueue.scala 150:36]
  wire [3:0] _GEN_871 = EntryValid_0 ? _GEN_755 : _GEN_188; // @[LoadStoreQueue.scala 150:36]
  wire [3:0] _GEN_872 = EntryValid_0 ? _GEN_756 : _GEN_189; // @[LoadStoreQueue.scala 150:36]
  wire [3:0] _GEN_873 = EntryValid_0 ? _GEN_757 : _GEN_190; // @[LoadStoreQueue.scala 150:36]
  wire [3:0] _GEN_874 = EntryValid_0 ? _GEN_758 : _GEN_191; // @[LoadStoreQueue.scala 150:36]
  wire [63:0] _GEN_875 = EntryValid_0 ? _GEN_759 : _GEN_218; // @[LoadStoreQueue.scala 150:36]
  wire [63:0] _GEN_876 = EntryValid_0 ? _GEN_760 : _GEN_230; // @[LoadStoreQueue.scala 150:36]
  wire [63:0] _GEN_877 = EntryValid_0 ? _GEN_761 : _GEN_242; // @[LoadStoreQueue.scala 150:36]
  wire [63:0] _GEN_878 = EntryValid_0 ? _GEN_762 : _GEN_254; // @[LoadStoreQueue.scala 150:36]
  wire [63:0] _GEN_879 = EntryValid_0 ? _GEN_763 : _GEN_266; // @[LoadStoreQueue.scala 150:36]
  wire [63:0] _GEN_880 = EntryValid_0 ? _GEN_764 : _GEN_278; // @[LoadStoreQueue.scala 150:36]
  wire [63:0] _GEN_881 = EntryValid_0 ? _GEN_765 : _GEN_290; // @[LoadStoreQueue.scala 150:36]
  wire [63:0] _GEN_882 = EntryValid_0 ? _GEN_766 : _GEN_302; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_883 = EntryValid_0 ? _GEN_767 : _GEN_219; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_884 = EntryValid_0 ? _GEN_768 : _GEN_231; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_885 = EntryValid_0 ? _GEN_769 : _GEN_243; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_886 = EntryValid_0 ? _GEN_770 : _GEN_255; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_887 = EntryValid_0 ? _GEN_771 : _GEN_267; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_888 = EntryValid_0 ? _GEN_772 : _GEN_279; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_889 = EntryValid_0 ? _GEN_773 : _GEN_291; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_890 = EntryValid_0 ? _GEN_774 : _GEN_303; // @[LoadStoreQueue.scala 150:36]
  wire [2:0] checkIndex_1 = nextTail + 3'h1; // @[LoadStoreQueue.scala 148:27]
  wire  _GEN_892 = 3'h1 == checkIndex_1 ? buffer_1_valid : buffer_0_valid; // @[LoadStoreQueue.scala 150:{36,36}]
  wire  _GEN_893 = 3'h2 == checkIndex_1 ? buffer_2_valid : _GEN_892; // @[LoadStoreQueue.scala 150:{36,36}]
  wire  _GEN_894 = 3'h3 == checkIndex_1 ? buffer_3_valid : _GEN_893; // @[LoadStoreQueue.scala 150:{36,36}]
  wire  _GEN_895 = 3'h4 == checkIndex_1 ? buffer_4_valid : _GEN_894; // @[LoadStoreQueue.scala 150:{36,36}]
  wire  _GEN_896 = 3'h5 == checkIndex_1 ? buffer_5_valid : _GEN_895; // @[LoadStoreQueue.scala 150:{36,36}]
  wire  _GEN_897 = 3'h6 == checkIndex_1 ? buffer_6_valid : _GEN_896; // @[LoadStoreQueue.scala 150:{36,36}]
  wire  EntryValid_1 = 3'h7 == checkIndex_1 ? buffer_7_valid : _GEN_897; // @[LoadStoreQueue.scala 150:{36,36}]
  wire [63:0] _GEN_900 = 3'h1 == checkIndex_1 ? buffer_1_address : buffer_0_address; // @[LoadStoreQueue.scala 151:{18,18}]
  wire [63:0] _GEN_901 = 3'h2 == checkIndex_1 ? buffer_2_address : _GEN_900; // @[LoadStoreQueue.scala 151:{18,18}]
  wire [63:0] _GEN_902 = 3'h3 == checkIndex_1 ? buffer_3_address : _GEN_901; // @[LoadStoreQueue.scala 151:{18,18}]
  wire [63:0] _GEN_903 = 3'h4 == checkIndex_1 ? buffer_4_address : _GEN_902; // @[LoadStoreQueue.scala 151:{18,18}]
  wire [63:0] _GEN_904 = 3'h5 == checkIndex_1 ? buffer_5_address : _GEN_903; // @[LoadStoreQueue.scala 151:{18,18}]
  wire [63:0] _GEN_905 = 3'h6 == checkIndex_1 ? buffer_6_address : _GEN_904; // @[LoadStoreQueue.scala 151:{18,18}]
  wire [63:0] _GEN_906 = 3'h7 == checkIndex_1 ? buffer_7_address : _GEN_905; // @[LoadStoreQueue.scala 151:{18,18}]
  wire  _GEN_908 = 3'h1 == checkIndex_1 ? buffer_1_addressValid : buffer_0_addressValid; // @[LoadStoreQueue.scala 152:{23,23}]
  wire  _GEN_909 = 3'h2 == checkIndex_1 ? buffer_2_addressValid : _GEN_908; // @[LoadStoreQueue.scala 152:{23,23}]
  wire  _GEN_910 = 3'h3 == checkIndex_1 ? buffer_3_addressValid : _GEN_909; // @[LoadStoreQueue.scala 152:{23,23}]
  wire  _GEN_911 = 3'h4 == checkIndex_1 ? buffer_4_addressValid : _GEN_910; // @[LoadStoreQueue.scala 152:{23,23}]
  wire  _GEN_912 = 3'h5 == checkIndex_1 ? buffer_5_addressValid : _GEN_911; // @[LoadStoreQueue.scala 152:{23,23}]
  wire  _GEN_913 = 3'h6 == checkIndex_1 ? buffer_6_addressValid : _GEN_912; // @[LoadStoreQueue.scala 152:{23,23}]
  wire  _GEN_914 = 3'h7 == checkIndex_1 ? buffer_7_addressValid : _GEN_913; // @[LoadStoreQueue.scala 152:{23,23}]
  wire  _T_237 = AddressValid_0 & Address_0 == _GEN_906; // @[LoadStoreQueue.scala 160:32]
  wire  _T_239 = _T_237 | ~AddressValid_0; // @[LoadStoreQueue.scala 162:26]
  wire  _GEN_916 = EntryValid_0 & _T_239; // @[LoadStoreQueue.scala 127:25 158:31]
  wire  _checkOk_T_13 = head != nextTail & EntryValid_1 & _GEN_914; // @[LoadStoreQueue.scala 171:62]
  wire  _GEN_918 = 3'h1 == checkIndex_1 ? buffer_1_info_accessType : buffer_0_info_accessType; // @[LoadStoreQueue.scala 174:{46,46}]
  wire  _GEN_919 = 3'h2 == checkIndex_1 ? buffer_2_info_accessType : _GEN_918; // @[LoadStoreQueue.scala 174:{46,46}]
  wire  _GEN_920 = 3'h3 == checkIndex_1 ? buffer_3_info_accessType : _GEN_919; // @[LoadStoreQueue.scala 174:{46,46}]
  wire  _GEN_921 = 3'h4 == checkIndex_1 ? buffer_4_info_accessType : _GEN_920; // @[LoadStoreQueue.scala 174:{46,46}]
  wire  _GEN_922 = 3'h5 == checkIndex_1 ? buffer_5_info_accessType : _GEN_921; // @[LoadStoreQueue.scala 174:{46,46}]
  wire  _GEN_923 = 3'h6 == checkIndex_1 ? buffer_6_info_accessType : _GEN_922; // @[LoadStoreQueue.scala 174:{46,46}]
  wire  _GEN_924 = 3'h7 == checkIndex_1 ? buffer_7_info_accessType : _GEN_923; // @[LoadStoreQueue.scala 174:{46,46}]
  wire  Overlap_1 = EntryValid_1 & _GEN_916; // @[LoadStoreQueue.scala 127:25 150:36]
  wire  _GEN_926 = 3'h1 == checkIndex_1 ? buffer_1_storeDataValid : buffer_0_storeDataValid; // @[LoadStoreQueue.scala 175:{57,57}]
  wire  _GEN_927 = 3'h2 == checkIndex_1 ? buffer_2_storeDataValid : _GEN_926; // @[LoadStoreQueue.scala 175:{57,57}]
  wire  _GEN_928 = 3'h3 == checkIndex_1 ? buffer_3_storeDataValid : _GEN_927; // @[LoadStoreQueue.scala 175:{57,57}]
  wire  _GEN_929 = 3'h4 == checkIndex_1 ? buffer_4_storeDataValid : _GEN_928; // @[LoadStoreQueue.scala 175:{57,57}]
  wire  _GEN_930 = 3'h5 == checkIndex_1 ? buffer_5_storeDataValid : _GEN_929; // @[LoadStoreQueue.scala 175:{57,57}]
  wire  _GEN_931 = 3'h6 == checkIndex_1 ? buffer_6_storeDataValid : _GEN_930; // @[LoadStoreQueue.scala 175:{57,57}]
  wire  _GEN_932 = 3'h7 == checkIndex_1 ? buffer_7_storeDataValid : _GEN_931; // @[LoadStoreQueue.scala 175:{57,57}]
  wire  _checkOk_T_18 = ~_GEN_924 & _GEN_932; // @[LoadStoreQueue.scala 175:57]
  wire  _GEN_934 = 3'h1 == checkIndex_1 ? buffer_1_readyReorderSign : buffer_0_readyReorderSign; // @[LoadStoreQueue.scala 177:{28,28}]
  wire  _GEN_935 = 3'h2 == checkIndex_1 ? buffer_2_readyReorderSign : _GEN_934; // @[LoadStoreQueue.scala 177:{28,28}]
  wire  _GEN_936 = 3'h3 == checkIndex_1 ? buffer_3_readyReorderSign : _GEN_935; // @[LoadStoreQueue.scala 177:{28,28}]
  wire  _GEN_937 = 3'h4 == checkIndex_1 ? buffer_4_readyReorderSign : _GEN_936; // @[LoadStoreQueue.scala 177:{28,28}]
  wire  _GEN_938 = 3'h5 == checkIndex_1 ? buffer_5_readyReorderSign : _GEN_937; // @[LoadStoreQueue.scala 177:{28,28}]
  wire  _GEN_939 = 3'h6 == checkIndex_1 ? buffer_6_readyReorderSign : _GEN_938; // @[LoadStoreQueue.scala 177:{28,28}]
  wire  _GEN_940 = 3'h7 == checkIndex_1 ? buffer_7_readyReorderSign : _GEN_939; // @[LoadStoreQueue.scala 177:{28,28}]
  wire  _checkOk_T_19 = _checkOk_T_18 & _GEN_940; // @[LoadStoreQueue.scala 177:28]
  wire  _checkOk_T_20 = _GEN_924 & ~Overlap_1 | _checkOk_T_19; // @[LoadStoreQueue.scala 174:71]
  wire  _checkOk_T_21 = _checkOk_T_13 & _checkOk_T_20; // @[LoadStoreQueue.scala 173:22]
  wire  checkOk_1 = EntryValid_1 & _checkOk_T_21; // @[LoadStoreQueue.scala 150:36 171:15 149:30]
  wire  _GEN_942 = 3'h1 == checkIndex_1 ? buffer_1_addressAndLoadResultTag_threadId :
    buffer_0_addressAndLoadResultTag_threadId; // @[LoadStoreQueue.scala 182:{28,28}]
  wire  _GEN_943 = 3'h2 == checkIndex_1 ? buffer_2_addressAndLoadResultTag_threadId : _GEN_942; // @[LoadStoreQueue.scala 182:{28,28}]
  wire  _GEN_944 = 3'h3 == checkIndex_1 ? buffer_3_addressAndLoadResultTag_threadId : _GEN_943; // @[LoadStoreQueue.scala 182:{28,28}]
  wire  _GEN_945 = 3'h4 == checkIndex_1 ? buffer_4_addressAndLoadResultTag_threadId : _GEN_944; // @[LoadStoreQueue.scala 182:{28,28}]
  wire  _GEN_946 = 3'h5 == checkIndex_1 ? buffer_5_addressAndLoadResultTag_threadId : _GEN_945; // @[LoadStoreQueue.scala 182:{28,28}]
  wire  _GEN_947 = 3'h6 == checkIndex_1 ? buffer_6_addressAndLoadResultTag_threadId : _GEN_946; // @[LoadStoreQueue.scala 182:{28,28}]
  wire  _GEN_948 = 3'h7 == checkIndex_1 ? buffer_7_addressAndLoadResultTag_threadId : _GEN_947; // @[LoadStoreQueue.scala 182:{28,28}]
  wire [3:0] _GEN_950 = 3'h1 == checkIndex_1 ? buffer_1_addressAndLoadResultTag_id : buffer_0_addressAndLoadResultTag_id
    ; // @[LoadStoreQueue.scala 182:{28,28}]
  wire [3:0] _GEN_951 = 3'h2 == checkIndex_1 ? buffer_2_addressAndLoadResultTag_id : _GEN_950; // @[LoadStoreQueue.scala 182:{28,28}]
  wire [3:0] _GEN_952 = 3'h3 == checkIndex_1 ? buffer_3_addressAndLoadResultTag_id : _GEN_951; // @[LoadStoreQueue.scala 182:{28,28}]
  wire [3:0] _GEN_953 = 3'h4 == checkIndex_1 ? buffer_4_addressAndLoadResultTag_id : _GEN_952; // @[LoadStoreQueue.scala 182:{28,28}]
  wire [3:0] _GEN_954 = 3'h5 == checkIndex_1 ? buffer_5_addressAndLoadResultTag_id : _GEN_953; // @[LoadStoreQueue.scala 182:{28,28}]
  wire [3:0] _GEN_955 = 3'h6 == checkIndex_1 ? buffer_6_addressAndLoadResultTag_id : _GEN_954; // @[LoadStoreQueue.scala 182:{28,28}]
  wire [3:0] _GEN_956 = 3'h7 == checkIndex_1 ? buffer_7_addressAndLoadResultTag_id : _GEN_955; // @[LoadStoreQueue.scala 182:{28,28}]
  wire [63:0] _GEN_958 = 3'h1 == checkIndex_1 ? buffer_1_storeData : buffer_0_storeData; // @[LoadStoreQueue.scala 183:{29,29}]
  wire [63:0] _GEN_959 = 3'h2 == checkIndex_1 ? buffer_2_storeData : _GEN_958; // @[LoadStoreQueue.scala 183:{29,29}]
  wire [63:0] _GEN_960 = 3'h3 == checkIndex_1 ? buffer_3_storeData : _GEN_959; // @[LoadStoreQueue.scala 183:{29,29}]
  wire [63:0] _GEN_961 = 3'h4 == checkIndex_1 ? buffer_4_storeData : _GEN_960; // @[LoadStoreQueue.scala 183:{29,29}]
  wire [63:0] _GEN_962 = 3'h5 == checkIndex_1 ? buffer_5_storeData : _GEN_961; // @[LoadStoreQueue.scala 183:{29,29}]
  wire [63:0] _GEN_963 = 3'h6 == checkIndex_1 ? buffer_6_storeData : _GEN_962; // @[LoadStoreQueue.scala 183:{29,29}]
  wire [63:0] _GEN_964 = 3'h7 == checkIndex_1 ? buffer_7_storeData : _GEN_963; // @[LoadStoreQueue.scala 183:{29,29}]
  wire  _GEN_966 = 3'h1 == checkIndex_1 ? buffer_1_info_signed : buffer_0_info_signed; // @[LoadStoreQueue.scala 185:{35,35}]
  wire  _GEN_967 = 3'h2 == checkIndex_1 ? buffer_2_info_signed : _GEN_966; // @[LoadStoreQueue.scala 185:{35,35}]
  wire  _GEN_968 = 3'h3 == checkIndex_1 ? buffer_3_info_signed : _GEN_967; // @[LoadStoreQueue.scala 185:{35,35}]
  wire  _GEN_969 = 3'h4 == checkIndex_1 ? buffer_4_info_signed : _GEN_968; // @[LoadStoreQueue.scala 185:{35,35}]
  wire  _GEN_970 = 3'h5 == checkIndex_1 ? buffer_5_info_signed : _GEN_969; // @[LoadStoreQueue.scala 185:{35,35}]
  wire  _GEN_971 = 3'h6 == checkIndex_1 ? buffer_6_info_signed : _GEN_970; // @[LoadStoreQueue.scala 185:{35,35}]
  wire  _GEN_972 = 3'h7 == checkIndex_1 ? buffer_7_info_signed : _GEN_971; // @[LoadStoreQueue.scala 185:{35,35}]
  wire [1:0] _GEN_974 = 3'h1 == checkIndex_1 ? buffer_1_info_accessWidth : buffer_0_info_accessWidth; // @[LoadStoreQueue.scala 185:{35,35}]
  wire [1:0] _GEN_975 = 3'h2 == checkIndex_1 ? buffer_2_info_accessWidth : _GEN_974; // @[LoadStoreQueue.scala 185:{35,35}]
  wire [1:0] _GEN_976 = 3'h3 == checkIndex_1 ? buffer_3_info_accessWidth : _GEN_975; // @[LoadStoreQueue.scala 185:{35,35}]
  wire [1:0] _GEN_977 = 3'h4 == checkIndex_1 ? buffer_4_info_accessWidth : _GEN_976; // @[LoadStoreQueue.scala 185:{35,35}]
  wire [1:0] _GEN_978 = 3'h5 == checkIndex_1 ? buffer_5_info_accessWidth : _GEN_977; // @[LoadStoreQueue.scala 185:{35,35}]
  wire [1:0] _GEN_979 = 3'h6 == checkIndex_1 ? buffer_6_info_accessWidth : _GEN_978; // @[LoadStoreQueue.scala 185:{35,35}]
  wire [1:0] _GEN_980 = 3'h7 == checkIndex_1 ? buffer_7_info_accessWidth : _GEN_979; // @[LoadStoreQueue.scala 185:{35,35}]
  wire  _GEN_981 = 3'h0 == checkIndex_1 ? 1'h0 : _GEN_787; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_982 = 3'h1 == checkIndex_1 ? 1'h0 : _GEN_788; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_983 = 3'h2 == checkIndex_1 ? 1'h0 : _GEN_789; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_984 = 3'h3 == checkIndex_1 ? 1'h0 : _GEN_790; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_985 = 3'h4 == checkIndex_1 ? 1'h0 : _GEN_791; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_986 = 3'h5 == checkIndex_1 ? 1'h0 : _GEN_792; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_987 = 3'h6 == checkIndex_1 ? 1'h0 : _GEN_793; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_988 = 3'h7 == checkIndex_1 ? 1'h0 : _GEN_794; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_989 = 3'h0 == checkIndex_1 ? 1'h0 : _GEN_795; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_990 = 3'h1 == checkIndex_1 ? 1'h0 : _GEN_796; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_991 = 3'h2 == checkIndex_1 ? 1'h0 : _GEN_797; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_992 = 3'h3 == checkIndex_1 ? 1'h0 : _GEN_798; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_993 = 3'h4 == checkIndex_1 ? 1'h0 : _GEN_799; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_994 = 3'h5 == checkIndex_1 ? 1'h0 : _GEN_800; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_995 = 3'h6 == checkIndex_1 ? 1'h0 : _GEN_801; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_996 = 3'h7 == checkIndex_1 ? 1'h0 : _GEN_802; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_997 = 3'h0 == checkIndex_1 ? 1'h0 : _GEN_803; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_998 = 3'h1 == checkIndex_1 ? 1'h0 : _GEN_804; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_999 = 3'h2 == checkIndex_1 ? 1'h0 : _GEN_805; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1000 = 3'h3 == checkIndex_1 ? 1'h0 : _GEN_806; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1001 = 3'h4 == checkIndex_1 ? 1'h0 : _GEN_807; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1002 = 3'h5 == checkIndex_1 ? 1'h0 : _GEN_808; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1003 = 3'h6 == checkIndex_1 ? 1'h0 : _GEN_809; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1004 = 3'h7 == checkIndex_1 ? 1'h0 : _GEN_810; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1005 = 3'h0 == checkIndex_1 ? 1'h0 : _GEN_811; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1006 = 3'h1 == checkIndex_1 ? 1'h0 : _GEN_812; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1007 = 3'h2 == checkIndex_1 ? 1'h0 : _GEN_813; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1008 = 3'h3 == checkIndex_1 ? 1'h0 : _GEN_814; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1009 = 3'h4 == checkIndex_1 ? 1'h0 : _GEN_815; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1010 = 3'h5 == checkIndex_1 ? 1'h0 : _GEN_816; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1011 = 3'h6 == checkIndex_1 ? 1'h0 : _GEN_817; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1012 = 3'h7 == checkIndex_1 ? 1'h0 : _GEN_818; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [1:0] _GEN_1013 = 3'h0 == checkIndex_1 ? 2'h0 : _GEN_819; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [1:0] _GEN_1014 = 3'h1 == checkIndex_1 ? 2'h0 : _GEN_820; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [1:0] _GEN_1015 = 3'h2 == checkIndex_1 ? 2'h0 : _GEN_821; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [1:0] _GEN_1016 = 3'h3 == checkIndex_1 ? 2'h0 : _GEN_822; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [1:0] _GEN_1017 = 3'h4 == checkIndex_1 ? 2'h0 : _GEN_823; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [1:0] _GEN_1018 = 3'h5 == checkIndex_1 ? 2'h0 : _GEN_824; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [1:0] _GEN_1019 = 3'h6 == checkIndex_1 ? 2'h0 : _GEN_825; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [1:0] _GEN_1020 = 3'h7 == checkIndex_1 ? 2'h0 : _GEN_826; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1021 = 3'h0 == checkIndex_1 ? 1'h0 : _GEN_827; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1022 = 3'h1 == checkIndex_1 ? 1'h0 : _GEN_828; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1023 = 3'h2 == checkIndex_1 ? 1'h0 : _GEN_829; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1024 = 3'h3 == checkIndex_1 ? 1'h0 : _GEN_830; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1025 = 3'h4 == checkIndex_1 ? 1'h0 : _GEN_831; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1026 = 3'h5 == checkIndex_1 ? 1'h0 : _GEN_832; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1027 = 3'h6 == checkIndex_1 ? 1'h0 : _GEN_833; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1028 = 3'h7 == checkIndex_1 ? 1'h0 : _GEN_834; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [3:0] _GEN_1029 = 3'h0 == checkIndex_1 ? 4'h0 : _GEN_835; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [3:0] _GEN_1030 = 3'h1 == checkIndex_1 ? 4'h0 : _GEN_836; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [3:0] _GEN_1031 = 3'h2 == checkIndex_1 ? 4'h0 : _GEN_837; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [3:0] _GEN_1032 = 3'h3 == checkIndex_1 ? 4'h0 : _GEN_838; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [3:0] _GEN_1033 = 3'h4 == checkIndex_1 ? 4'h0 : _GEN_839; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [3:0] _GEN_1034 = 3'h5 == checkIndex_1 ? 4'h0 : _GEN_840; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [3:0] _GEN_1035 = 3'h6 == checkIndex_1 ? 4'h0 : _GEN_841; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [3:0] _GEN_1036 = 3'h7 == checkIndex_1 ? 4'h0 : _GEN_842; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [63:0] _GEN_1037 = 3'h0 == checkIndex_1 ? 64'h0 : _GEN_843; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [63:0] _GEN_1038 = 3'h1 == checkIndex_1 ? 64'h0 : _GEN_844; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [63:0] _GEN_1039 = 3'h2 == checkIndex_1 ? 64'h0 : _GEN_845; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [63:0] _GEN_1040 = 3'h3 == checkIndex_1 ? 64'h0 : _GEN_846; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [63:0] _GEN_1041 = 3'h4 == checkIndex_1 ? 64'h0 : _GEN_847; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [63:0] _GEN_1042 = 3'h5 == checkIndex_1 ? 64'h0 : _GEN_848; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [63:0] _GEN_1043 = 3'h6 == checkIndex_1 ? 64'h0 : _GEN_849; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [63:0] _GEN_1044 = 3'h7 == checkIndex_1 ? 64'h0 : _GEN_850; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1045 = 3'h0 == checkIndex_1 ? 1'h0 : _GEN_851; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1046 = 3'h1 == checkIndex_1 ? 1'h0 : _GEN_852; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1047 = 3'h2 == checkIndex_1 ? 1'h0 : _GEN_853; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1048 = 3'h3 == checkIndex_1 ? 1'h0 : _GEN_854; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1049 = 3'h4 == checkIndex_1 ? 1'h0 : _GEN_855; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1050 = 3'h5 == checkIndex_1 ? 1'h0 : _GEN_856; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1051 = 3'h6 == checkIndex_1 ? 1'h0 : _GEN_857; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1052 = 3'h7 == checkIndex_1 ? 1'h0 : _GEN_858; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1053 = 3'h0 == checkIndex_1 ? 1'h0 : _GEN_859; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1054 = 3'h1 == checkIndex_1 ? 1'h0 : _GEN_860; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1055 = 3'h2 == checkIndex_1 ? 1'h0 : _GEN_861; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1056 = 3'h3 == checkIndex_1 ? 1'h0 : _GEN_862; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1057 = 3'h4 == checkIndex_1 ? 1'h0 : _GEN_863; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1058 = 3'h5 == checkIndex_1 ? 1'h0 : _GEN_864; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1059 = 3'h6 == checkIndex_1 ? 1'h0 : _GEN_865; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1060 = 3'h7 == checkIndex_1 ? 1'h0 : _GEN_866; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [3:0] _GEN_1061 = 3'h0 == checkIndex_1 ? 4'h0 : _GEN_867; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [3:0] _GEN_1062 = 3'h1 == checkIndex_1 ? 4'h0 : _GEN_868; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [3:0] _GEN_1063 = 3'h2 == checkIndex_1 ? 4'h0 : _GEN_869; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [3:0] _GEN_1064 = 3'h3 == checkIndex_1 ? 4'h0 : _GEN_870; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [3:0] _GEN_1065 = 3'h4 == checkIndex_1 ? 4'h0 : _GEN_871; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [3:0] _GEN_1066 = 3'h5 == checkIndex_1 ? 4'h0 : _GEN_872; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [3:0] _GEN_1067 = 3'h6 == checkIndex_1 ? 4'h0 : _GEN_873; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [3:0] _GEN_1068 = 3'h7 == checkIndex_1 ? 4'h0 : _GEN_874; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [63:0] _GEN_1069 = 3'h0 == checkIndex_1 ? 64'h0 : _GEN_875; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [63:0] _GEN_1070 = 3'h1 == checkIndex_1 ? 64'h0 : _GEN_876; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [63:0] _GEN_1071 = 3'h2 == checkIndex_1 ? 64'h0 : _GEN_877; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [63:0] _GEN_1072 = 3'h3 == checkIndex_1 ? 64'h0 : _GEN_878; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [63:0] _GEN_1073 = 3'h4 == checkIndex_1 ? 64'h0 : _GEN_879; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [63:0] _GEN_1074 = 3'h5 == checkIndex_1 ? 64'h0 : _GEN_880; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [63:0] _GEN_1075 = 3'h6 == checkIndex_1 ? 64'h0 : _GEN_881; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [63:0] _GEN_1076 = 3'h7 == checkIndex_1 ? 64'h0 : _GEN_882; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1077 = 3'h0 == checkIndex_1 ? 1'h0 : _GEN_883; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1078 = 3'h1 == checkIndex_1 ? 1'h0 : _GEN_884; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1079 = 3'h2 == checkIndex_1 ? 1'h0 : _GEN_885; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1080 = 3'h3 == checkIndex_1 ? 1'h0 : _GEN_886; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1081 = 3'h4 == checkIndex_1 ? 1'h0 : _GEN_887; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1082 = 3'h5 == checkIndex_1 ? 1'h0 : _GEN_888; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1083 = 3'h6 == checkIndex_1 ? 1'h0 : _GEN_889; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1084 = 3'h7 == checkIndex_1 ? 1'h0 : _GEN_890; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1085 = io_memory_ready ? _GEN_981 : _GEN_787; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_1086 = io_memory_ready ? _GEN_982 : _GEN_788; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_1087 = io_memory_ready ? _GEN_983 : _GEN_789; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_1088 = io_memory_ready ? _GEN_984 : _GEN_790; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_1089 = io_memory_ready ? _GEN_985 : _GEN_791; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_1090 = io_memory_ready ? _GEN_986 : _GEN_792; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_1091 = io_memory_ready ? _GEN_987 : _GEN_793; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_1092 = io_memory_ready ? _GEN_988 : _GEN_794; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_1093 = io_memory_ready ? _GEN_989 : _GEN_795; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_1094 = io_memory_ready ? _GEN_990 : _GEN_796; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_1095 = io_memory_ready ? _GEN_991 : _GEN_797; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_1096 = io_memory_ready ? _GEN_992 : _GEN_798; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_1097 = io_memory_ready ? _GEN_993 : _GEN_799; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_1098 = io_memory_ready ? _GEN_994 : _GEN_800; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_1099 = io_memory_ready ? _GEN_995 : _GEN_801; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_1100 = io_memory_ready ? _GEN_996 : _GEN_802; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_1101 = io_memory_ready ? _GEN_997 : _GEN_803; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_1102 = io_memory_ready ? _GEN_998 : _GEN_804; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_1103 = io_memory_ready ? _GEN_999 : _GEN_805; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_1104 = io_memory_ready ? _GEN_1000 : _GEN_806; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_1105 = io_memory_ready ? _GEN_1001 : _GEN_807; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_1106 = io_memory_ready ? _GEN_1002 : _GEN_808; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_1107 = io_memory_ready ? _GEN_1003 : _GEN_809; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_1108 = io_memory_ready ? _GEN_1004 : _GEN_810; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_1109 = io_memory_ready ? _GEN_1005 : _GEN_811; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_1110 = io_memory_ready ? _GEN_1006 : _GEN_812; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_1111 = io_memory_ready ? _GEN_1007 : _GEN_813; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_1112 = io_memory_ready ? _GEN_1008 : _GEN_814; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_1113 = io_memory_ready ? _GEN_1009 : _GEN_815; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_1114 = io_memory_ready ? _GEN_1010 : _GEN_816; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_1115 = io_memory_ready ? _GEN_1011 : _GEN_817; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_1116 = io_memory_ready ? _GEN_1012 : _GEN_818; // @[LoadStoreQueue.scala 186:31]
  wire [1:0] _GEN_1117 = io_memory_ready ? _GEN_1013 : _GEN_819; // @[LoadStoreQueue.scala 186:31]
  wire [1:0] _GEN_1118 = io_memory_ready ? _GEN_1014 : _GEN_820; // @[LoadStoreQueue.scala 186:31]
  wire [1:0] _GEN_1119 = io_memory_ready ? _GEN_1015 : _GEN_821; // @[LoadStoreQueue.scala 186:31]
  wire [1:0] _GEN_1120 = io_memory_ready ? _GEN_1016 : _GEN_822; // @[LoadStoreQueue.scala 186:31]
  wire [1:0] _GEN_1121 = io_memory_ready ? _GEN_1017 : _GEN_823; // @[LoadStoreQueue.scala 186:31]
  wire [1:0] _GEN_1122 = io_memory_ready ? _GEN_1018 : _GEN_824; // @[LoadStoreQueue.scala 186:31]
  wire [1:0] _GEN_1123 = io_memory_ready ? _GEN_1019 : _GEN_825; // @[LoadStoreQueue.scala 186:31]
  wire [1:0] _GEN_1124 = io_memory_ready ? _GEN_1020 : _GEN_826; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_1125 = io_memory_ready ? _GEN_1021 : _GEN_827; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_1126 = io_memory_ready ? _GEN_1022 : _GEN_828; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_1127 = io_memory_ready ? _GEN_1023 : _GEN_829; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_1128 = io_memory_ready ? _GEN_1024 : _GEN_830; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_1129 = io_memory_ready ? _GEN_1025 : _GEN_831; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_1130 = io_memory_ready ? _GEN_1026 : _GEN_832; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_1131 = io_memory_ready ? _GEN_1027 : _GEN_833; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_1132 = io_memory_ready ? _GEN_1028 : _GEN_834; // @[LoadStoreQueue.scala 186:31]
  wire [3:0] _GEN_1133 = io_memory_ready ? _GEN_1029 : _GEN_835; // @[LoadStoreQueue.scala 186:31]
  wire [3:0] _GEN_1134 = io_memory_ready ? _GEN_1030 : _GEN_836; // @[LoadStoreQueue.scala 186:31]
  wire [3:0] _GEN_1135 = io_memory_ready ? _GEN_1031 : _GEN_837; // @[LoadStoreQueue.scala 186:31]
  wire [3:0] _GEN_1136 = io_memory_ready ? _GEN_1032 : _GEN_838; // @[LoadStoreQueue.scala 186:31]
  wire [3:0] _GEN_1137 = io_memory_ready ? _GEN_1033 : _GEN_839; // @[LoadStoreQueue.scala 186:31]
  wire [3:0] _GEN_1138 = io_memory_ready ? _GEN_1034 : _GEN_840; // @[LoadStoreQueue.scala 186:31]
  wire [3:0] _GEN_1139 = io_memory_ready ? _GEN_1035 : _GEN_841; // @[LoadStoreQueue.scala 186:31]
  wire [3:0] _GEN_1140 = io_memory_ready ? _GEN_1036 : _GEN_842; // @[LoadStoreQueue.scala 186:31]
  wire [63:0] _GEN_1141 = io_memory_ready ? _GEN_1037 : _GEN_843; // @[LoadStoreQueue.scala 186:31]
  wire [63:0] _GEN_1142 = io_memory_ready ? _GEN_1038 : _GEN_844; // @[LoadStoreQueue.scala 186:31]
  wire [63:0] _GEN_1143 = io_memory_ready ? _GEN_1039 : _GEN_845; // @[LoadStoreQueue.scala 186:31]
  wire [63:0] _GEN_1144 = io_memory_ready ? _GEN_1040 : _GEN_846; // @[LoadStoreQueue.scala 186:31]
  wire [63:0] _GEN_1145 = io_memory_ready ? _GEN_1041 : _GEN_847; // @[LoadStoreQueue.scala 186:31]
  wire [63:0] _GEN_1146 = io_memory_ready ? _GEN_1042 : _GEN_848; // @[LoadStoreQueue.scala 186:31]
  wire [63:0] _GEN_1147 = io_memory_ready ? _GEN_1043 : _GEN_849; // @[LoadStoreQueue.scala 186:31]
  wire [63:0] _GEN_1148 = io_memory_ready ? _GEN_1044 : _GEN_850; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_1149 = io_memory_ready ? _GEN_1045 : _GEN_851; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_1150 = io_memory_ready ? _GEN_1046 : _GEN_852; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_1151 = io_memory_ready ? _GEN_1047 : _GEN_853; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_1152 = io_memory_ready ? _GEN_1048 : _GEN_854; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_1153 = io_memory_ready ? _GEN_1049 : _GEN_855; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_1154 = io_memory_ready ? _GEN_1050 : _GEN_856; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_1155 = io_memory_ready ? _GEN_1051 : _GEN_857; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_1156 = io_memory_ready ? _GEN_1052 : _GEN_858; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_1157 = io_memory_ready ? _GEN_1053 : _GEN_859; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_1158 = io_memory_ready ? _GEN_1054 : _GEN_860; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_1159 = io_memory_ready ? _GEN_1055 : _GEN_861; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_1160 = io_memory_ready ? _GEN_1056 : _GEN_862; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_1161 = io_memory_ready ? _GEN_1057 : _GEN_863; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_1162 = io_memory_ready ? _GEN_1058 : _GEN_864; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_1163 = io_memory_ready ? _GEN_1059 : _GEN_865; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_1164 = io_memory_ready ? _GEN_1060 : _GEN_866; // @[LoadStoreQueue.scala 186:31]
  wire [3:0] _GEN_1165 = io_memory_ready ? _GEN_1061 : _GEN_867; // @[LoadStoreQueue.scala 186:31]
  wire [3:0] _GEN_1166 = io_memory_ready ? _GEN_1062 : _GEN_868; // @[LoadStoreQueue.scala 186:31]
  wire [3:0] _GEN_1167 = io_memory_ready ? _GEN_1063 : _GEN_869; // @[LoadStoreQueue.scala 186:31]
  wire [3:0] _GEN_1168 = io_memory_ready ? _GEN_1064 : _GEN_870; // @[LoadStoreQueue.scala 186:31]
  wire [3:0] _GEN_1169 = io_memory_ready ? _GEN_1065 : _GEN_871; // @[LoadStoreQueue.scala 186:31]
  wire [3:0] _GEN_1170 = io_memory_ready ? _GEN_1066 : _GEN_872; // @[LoadStoreQueue.scala 186:31]
  wire [3:0] _GEN_1171 = io_memory_ready ? _GEN_1067 : _GEN_873; // @[LoadStoreQueue.scala 186:31]
  wire [3:0] _GEN_1172 = io_memory_ready ? _GEN_1068 : _GEN_874; // @[LoadStoreQueue.scala 186:31]
  wire [63:0] _GEN_1173 = io_memory_ready ? _GEN_1069 : _GEN_875; // @[LoadStoreQueue.scala 186:31]
  wire [63:0] _GEN_1174 = io_memory_ready ? _GEN_1070 : _GEN_876; // @[LoadStoreQueue.scala 186:31]
  wire [63:0] _GEN_1175 = io_memory_ready ? _GEN_1071 : _GEN_877; // @[LoadStoreQueue.scala 186:31]
  wire [63:0] _GEN_1176 = io_memory_ready ? _GEN_1072 : _GEN_878; // @[LoadStoreQueue.scala 186:31]
  wire [63:0] _GEN_1177 = io_memory_ready ? _GEN_1073 : _GEN_879; // @[LoadStoreQueue.scala 186:31]
  wire [63:0] _GEN_1178 = io_memory_ready ? _GEN_1074 : _GEN_880; // @[LoadStoreQueue.scala 186:31]
  wire [63:0] _GEN_1179 = io_memory_ready ? _GEN_1075 : _GEN_881; // @[LoadStoreQueue.scala 186:31]
  wire [63:0] _GEN_1180 = io_memory_ready ? _GEN_1076 : _GEN_882; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_1181 = io_memory_ready ? _GEN_1077 : _GEN_883; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_1182 = io_memory_ready ? _GEN_1078 : _GEN_884; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_1183 = io_memory_ready ? _GEN_1079 : _GEN_885; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_1184 = io_memory_ready ? _GEN_1080 : _GEN_886; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_1185 = io_memory_ready ? _GEN_1081 : _GEN_887; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_1186 = io_memory_ready ? _GEN_1082 : _GEN_888; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_1187 = io_memory_ready ? _GEN_1083 : _GEN_889; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_1188 = io_memory_ready ? _GEN_1084 : _GEN_890; // @[LoadStoreQueue.scala 186:31]
  wire  _GEN_1189 = checkOk_1 & ~checkOk ? _GEN_948 : _GEN_423; // @[LoadStoreQueue.scala 181:31 182:28]
  wire [3:0] _GEN_1190 = checkOk_1 & ~checkOk ? _GEN_956 : _GEN_431; // @[LoadStoreQueue.scala 181:31 182:28]
  wire [63:0] _GEN_1191 = checkOk_1 & ~checkOk ? _GEN_964 : _GEN_439; // @[LoadStoreQueue.scala 181:31 183:29]
  wire [63:0] _GEN_1192 = checkOk_1 & ~checkOk ? _GEN_906 : _GEN_383; // @[LoadStoreQueue.scala 181:31 184:32]
  wire  _GEN_1193 = checkOk_1 & ~checkOk ? _GEN_924 : _GEN_399; // @[LoadStoreQueue.scala 181:31 185:35]
  wire  _GEN_1194 = checkOk_1 & ~checkOk ? _GEN_972 : _GEN_447; // @[LoadStoreQueue.scala 181:31 185:35]
  wire [1:0] _GEN_1195 = checkOk_1 & ~checkOk ? _GEN_980 : _GEN_455; // @[LoadStoreQueue.scala 181:31 185:35]
  wire  _GEN_1196 = checkOk_1 & ~checkOk ? _GEN_1085 : _GEN_787; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_1197 = checkOk_1 & ~checkOk ? _GEN_1086 : _GEN_788; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_1198 = checkOk_1 & ~checkOk ? _GEN_1087 : _GEN_789; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_1199 = checkOk_1 & ~checkOk ? _GEN_1088 : _GEN_790; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_1200 = checkOk_1 & ~checkOk ? _GEN_1089 : _GEN_791; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_1201 = checkOk_1 & ~checkOk ? _GEN_1090 : _GEN_792; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_1202 = checkOk_1 & ~checkOk ? _GEN_1091 : _GEN_793; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_1203 = checkOk_1 & ~checkOk ? _GEN_1092 : _GEN_794; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_1204 = checkOk_1 & ~checkOk ? _GEN_1093 : _GEN_795; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_1205 = checkOk_1 & ~checkOk ? _GEN_1094 : _GEN_796; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_1206 = checkOk_1 & ~checkOk ? _GEN_1095 : _GEN_797; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_1207 = checkOk_1 & ~checkOk ? _GEN_1096 : _GEN_798; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_1208 = checkOk_1 & ~checkOk ? _GEN_1097 : _GEN_799; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_1209 = checkOk_1 & ~checkOk ? _GEN_1098 : _GEN_800; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_1210 = checkOk_1 & ~checkOk ? _GEN_1099 : _GEN_801; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_1211 = checkOk_1 & ~checkOk ? _GEN_1100 : _GEN_802; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_1212 = checkOk_1 & ~checkOk ? _GEN_1101 : _GEN_803; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_1213 = checkOk_1 & ~checkOk ? _GEN_1102 : _GEN_804; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_1214 = checkOk_1 & ~checkOk ? _GEN_1103 : _GEN_805; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_1215 = checkOk_1 & ~checkOk ? _GEN_1104 : _GEN_806; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_1216 = checkOk_1 & ~checkOk ? _GEN_1105 : _GEN_807; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_1217 = checkOk_1 & ~checkOk ? _GEN_1106 : _GEN_808; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_1218 = checkOk_1 & ~checkOk ? _GEN_1107 : _GEN_809; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_1219 = checkOk_1 & ~checkOk ? _GEN_1108 : _GEN_810; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_1220 = checkOk_1 & ~checkOk ? _GEN_1109 : _GEN_811; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_1221 = checkOk_1 & ~checkOk ? _GEN_1110 : _GEN_812; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_1222 = checkOk_1 & ~checkOk ? _GEN_1111 : _GEN_813; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_1223 = checkOk_1 & ~checkOk ? _GEN_1112 : _GEN_814; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_1224 = checkOk_1 & ~checkOk ? _GEN_1113 : _GEN_815; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_1225 = checkOk_1 & ~checkOk ? _GEN_1114 : _GEN_816; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_1226 = checkOk_1 & ~checkOk ? _GEN_1115 : _GEN_817; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_1227 = checkOk_1 & ~checkOk ? _GEN_1116 : _GEN_818; // @[LoadStoreQueue.scala 181:31]
  wire [1:0] _GEN_1228 = checkOk_1 & ~checkOk ? _GEN_1117 : _GEN_819; // @[LoadStoreQueue.scala 181:31]
  wire [1:0] _GEN_1229 = checkOk_1 & ~checkOk ? _GEN_1118 : _GEN_820; // @[LoadStoreQueue.scala 181:31]
  wire [1:0] _GEN_1230 = checkOk_1 & ~checkOk ? _GEN_1119 : _GEN_821; // @[LoadStoreQueue.scala 181:31]
  wire [1:0] _GEN_1231 = checkOk_1 & ~checkOk ? _GEN_1120 : _GEN_822; // @[LoadStoreQueue.scala 181:31]
  wire [1:0] _GEN_1232 = checkOk_1 & ~checkOk ? _GEN_1121 : _GEN_823; // @[LoadStoreQueue.scala 181:31]
  wire [1:0] _GEN_1233 = checkOk_1 & ~checkOk ? _GEN_1122 : _GEN_824; // @[LoadStoreQueue.scala 181:31]
  wire [1:0] _GEN_1234 = checkOk_1 & ~checkOk ? _GEN_1123 : _GEN_825; // @[LoadStoreQueue.scala 181:31]
  wire [1:0] _GEN_1235 = checkOk_1 & ~checkOk ? _GEN_1124 : _GEN_826; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_1236 = checkOk_1 & ~checkOk ? _GEN_1125 : _GEN_827; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_1237 = checkOk_1 & ~checkOk ? _GEN_1126 : _GEN_828; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_1238 = checkOk_1 & ~checkOk ? _GEN_1127 : _GEN_829; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_1239 = checkOk_1 & ~checkOk ? _GEN_1128 : _GEN_830; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_1240 = checkOk_1 & ~checkOk ? _GEN_1129 : _GEN_831; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_1241 = checkOk_1 & ~checkOk ? _GEN_1130 : _GEN_832; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_1242 = checkOk_1 & ~checkOk ? _GEN_1131 : _GEN_833; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_1243 = checkOk_1 & ~checkOk ? _GEN_1132 : _GEN_834; // @[LoadStoreQueue.scala 181:31]
  wire [3:0] _GEN_1244 = checkOk_1 & ~checkOk ? _GEN_1133 : _GEN_835; // @[LoadStoreQueue.scala 181:31]
  wire [3:0] _GEN_1245 = checkOk_1 & ~checkOk ? _GEN_1134 : _GEN_836; // @[LoadStoreQueue.scala 181:31]
  wire [3:0] _GEN_1246 = checkOk_1 & ~checkOk ? _GEN_1135 : _GEN_837; // @[LoadStoreQueue.scala 181:31]
  wire [3:0] _GEN_1247 = checkOk_1 & ~checkOk ? _GEN_1136 : _GEN_838; // @[LoadStoreQueue.scala 181:31]
  wire [3:0] _GEN_1248 = checkOk_1 & ~checkOk ? _GEN_1137 : _GEN_839; // @[LoadStoreQueue.scala 181:31]
  wire [3:0] _GEN_1249 = checkOk_1 & ~checkOk ? _GEN_1138 : _GEN_840; // @[LoadStoreQueue.scala 181:31]
  wire [3:0] _GEN_1250 = checkOk_1 & ~checkOk ? _GEN_1139 : _GEN_841; // @[LoadStoreQueue.scala 181:31]
  wire [3:0] _GEN_1251 = checkOk_1 & ~checkOk ? _GEN_1140 : _GEN_842; // @[LoadStoreQueue.scala 181:31]
  wire [63:0] _GEN_1252 = checkOk_1 & ~checkOk ? _GEN_1141 : _GEN_843; // @[LoadStoreQueue.scala 181:31]
  wire [63:0] _GEN_1253 = checkOk_1 & ~checkOk ? _GEN_1142 : _GEN_844; // @[LoadStoreQueue.scala 181:31]
  wire [63:0] _GEN_1254 = checkOk_1 & ~checkOk ? _GEN_1143 : _GEN_845; // @[LoadStoreQueue.scala 181:31]
  wire [63:0] _GEN_1255 = checkOk_1 & ~checkOk ? _GEN_1144 : _GEN_846; // @[LoadStoreQueue.scala 181:31]
  wire [63:0] _GEN_1256 = checkOk_1 & ~checkOk ? _GEN_1145 : _GEN_847; // @[LoadStoreQueue.scala 181:31]
  wire [63:0] _GEN_1257 = checkOk_1 & ~checkOk ? _GEN_1146 : _GEN_848; // @[LoadStoreQueue.scala 181:31]
  wire [63:0] _GEN_1258 = checkOk_1 & ~checkOk ? _GEN_1147 : _GEN_849; // @[LoadStoreQueue.scala 181:31]
  wire [63:0] _GEN_1259 = checkOk_1 & ~checkOk ? _GEN_1148 : _GEN_850; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_1260 = checkOk_1 & ~checkOk ? _GEN_1149 : _GEN_851; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_1261 = checkOk_1 & ~checkOk ? _GEN_1150 : _GEN_852; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_1262 = checkOk_1 & ~checkOk ? _GEN_1151 : _GEN_853; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_1263 = checkOk_1 & ~checkOk ? _GEN_1152 : _GEN_854; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_1264 = checkOk_1 & ~checkOk ? _GEN_1153 : _GEN_855; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_1265 = checkOk_1 & ~checkOk ? _GEN_1154 : _GEN_856; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_1266 = checkOk_1 & ~checkOk ? _GEN_1155 : _GEN_857; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_1267 = checkOk_1 & ~checkOk ? _GEN_1156 : _GEN_858; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_1268 = checkOk_1 & ~checkOk ? _GEN_1157 : _GEN_859; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_1269 = checkOk_1 & ~checkOk ? _GEN_1158 : _GEN_860; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_1270 = checkOk_1 & ~checkOk ? _GEN_1159 : _GEN_861; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_1271 = checkOk_1 & ~checkOk ? _GEN_1160 : _GEN_862; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_1272 = checkOk_1 & ~checkOk ? _GEN_1161 : _GEN_863; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_1273 = checkOk_1 & ~checkOk ? _GEN_1162 : _GEN_864; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_1274 = checkOk_1 & ~checkOk ? _GEN_1163 : _GEN_865; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_1275 = checkOk_1 & ~checkOk ? _GEN_1164 : _GEN_866; // @[LoadStoreQueue.scala 181:31]
  wire [3:0] _GEN_1276 = checkOk_1 & ~checkOk ? _GEN_1165 : _GEN_867; // @[LoadStoreQueue.scala 181:31]
  wire [3:0] _GEN_1277 = checkOk_1 & ~checkOk ? _GEN_1166 : _GEN_868; // @[LoadStoreQueue.scala 181:31]
  wire [3:0] _GEN_1278 = checkOk_1 & ~checkOk ? _GEN_1167 : _GEN_869; // @[LoadStoreQueue.scala 181:31]
  wire [3:0] _GEN_1279 = checkOk_1 & ~checkOk ? _GEN_1168 : _GEN_870; // @[LoadStoreQueue.scala 181:31]
  wire [3:0] _GEN_1280 = checkOk_1 & ~checkOk ? _GEN_1169 : _GEN_871; // @[LoadStoreQueue.scala 181:31]
  wire [3:0] _GEN_1281 = checkOk_1 & ~checkOk ? _GEN_1170 : _GEN_872; // @[LoadStoreQueue.scala 181:31]
  wire [3:0] _GEN_1282 = checkOk_1 & ~checkOk ? _GEN_1171 : _GEN_873; // @[LoadStoreQueue.scala 181:31]
  wire [3:0] _GEN_1283 = checkOk_1 & ~checkOk ? _GEN_1172 : _GEN_874; // @[LoadStoreQueue.scala 181:31]
  wire [63:0] _GEN_1284 = checkOk_1 & ~checkOk ? _GEN_1173 : _GEN_875; // @[LoadStoreQueue.scala 181:31]
  wire [63:0] _GEN_1285 = checkOk_1 & ~checkOk ? _GEN_1174 : _GEN_876; // @[LoadStoreQueue.scala 181:31]
  wire [63:0] _GEN_1286 = checkOk_1 & ~checkOk ? _GEN_1175 : _GEN_877; // @[LoadStoreQueue.scala 181:31]
  wire [63:0] _GEN_1287 = checkOk_1 & ~checkOk ? _GEN_1176 : _GEN_878; // @[LoadStoreQueue.scala 181:31]
  wire [63:0] _GEN_1288 = checkOk_1 & ~checkOk ? _GEN_1177 : _GEN_879; // @[LoadStoreQueue.scala 181:31]
  wire [63:0] _GEN_1289 = checkOk_1 & ~checkOk ? _GEN_1178 : _GEN_880; // @[LoadStoreQueue.scala 181:31]
  wire [63:0] _GEN_1290 = checkOk_1 & ~checkOk ? _GEN_1179 : _GEN_881; // @[LoadStoreQueue.scala 181:31]
  wire [63:0] _GEN_1291 = checkOk_1 & ~checkOk ? _GEN_1180 : _GEN_882; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_1292 = checkOk_1 & ~checkOk ? _GEN_1181 : _GEN_883; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_1293 = checkOk_1 & ~checkOk ? _GEN_1182 : _GEN_884; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_1294 = checkOk_1 & ~checkOk ? _GEN_1183 : _GEN_885; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_1295 = checkOk_1 & ~checkOk ? _GEN_1184 : _GEN_886; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_1296 = checkOk_1 & ~checkOk ? _GEN_1185 : _GEN_887; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_1297 = checkOk_1 & ~checkOk ? _GEN_1186 : _GEN_888; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_1298 = checkOk_1 & ~checkOk ? _GEN_1187 : _GEN_889; // @[LoadStoreQueue.scala 181:31]
  wire  _GEN_1299 = checkOk_1 & ~checkOk ? _GEN_1188 : _GEN_890; // @[LoadStoreQueue.scala 181:31]
  wire [63:0] Address_1 = EntryValid_1 ? _GEN_906 : 64'h0; // @[LoadStoreQueue.scala 150:36 151:18 130:25]
  wire  AddressValid_1 = EntryValid_1 & _GEN_914; // @[LoadStoreQueue.scala 150:36 152:23 133:30]
  wire  _GEN_1305 = EntryValid_1 ? checkOk_1 | checkOk : _GEN_779; // @[LoadStoreQueue.scala 150:36 179:23]
  wire  _GEN_1306 = EntryValid_1 ? _GEN_1189 : _GEN_423; // @[LoadStoreQueue.scala 150:36]
  wire [3:0] _GEN_1307 = EntryValid_1 ? _GEN_1190 : _GEN_431; // @[LoadStoreQueue.scala 150:36]
  wire [63:0] _GEN_1308 = EntryValid_1 ? _GEN_1191 : _GEN_439; // @[LoadStoreQueue.scala 150:36]
  wire [63:0] _GEN_1309 = EntryValid_1 ? _GEN_1192 : _GEN_383; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1310 = EntryValid_1 ? _GEN_1193 : _GEN_399; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1311 = EntryValid_1 ? _GEN_1194 : _GEN_447; // @[LoadStoreQueue.scala 150:36]
  wire [1:0] _GEN_1312 = EntryValid_1 ? _GEN_1195 : _GEN_455; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1313 = EntryValid_1 ? _GEN_1196 : _GEN_787; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1314 = EntryValid_1 ? _GEN_1197 : _GEN_788; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1315 = EntryValid_1 ? _GEN_1198 : _GEN_789; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1316 = EntryValid_1 ? _GEN_1199 : _GEN_790; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1317 = EntryValid_1 ? _GEN_1200 : _GEN_791; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1318 = EntryValid_1 ? _GEN_1201 : _GEN_792; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1319 = EntryValid_1 ? _GEN_1202 : _GEN_793; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1320 = EntryValid_1 ? _GEN_1203 : _GEN_794; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1321 = EntryValid_1 ? _GEN_1204 : _GEN_795; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1322 = EntryValid_1 ? _GEN_1205 : _GEN_796; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1323 = EntryValid_1 ? _GEN_1206 : _GEN_797; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1324 = EntryValid_1 ? _GEN_1207 : _GEN_798; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1325 = EntryValid_1 ? _GEN_1208 : _GEN_799; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1326 = EntryValid_1 ? _GEN_1209 : _GEN_800; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1327 = EntryValid_1 ? _GEN_1210 : _GEN_801; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1328 = EntryValid_1 ? _GEN_1211 : _GEN_802; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1329 = EntryValid_1 ? _GEN_1212 : _GEN_803; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1330 = EntryValid_1 ? _GEN_1213 : _GEN_804; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1331 = EntryValid_1 ? _GEN_1214 : _GEN_805; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1332 = EntryValid_1 ? _GEN_1215 : _GEN_806; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1333 = EntryValid_1 ? _GEN_1216 : _GEN_807; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1334 = EntryValid_1 ? _GEN_1217 : _GEN_808; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1335 = EntryValid_1 ? _GEN_1218 : _GEN_809; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1336 = EntryValid_1 ? _GEN_1219 : _GEN_810; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1337 = EntryValid_1 ? _GEN_1220 : _GEN_811; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1338 = EntryValid_1 ? _GEN_1221 : _GEN_812; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1339 = EntryValid_1 ? _GEN_1222 : _GEN_813; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1340 = EntryValid_1 ? _GEN_1223 : _GEN_814; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1341 = EntryValid_1 ? _GEN_1224 : _GEN_815; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1342 = EntryValid_1 ? _GEN_1225 : _GEN_816; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1343 = EntryValid_1 ? _GEN_1226 : _GEN_817; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1344 = EntryValid_1 ? _GEN_1227 : _GEN_818; // @[LoadStoreQueue.scala 150:36]
  wire [1:0] _GEN_1345 = EntryValid_1 ? _GEN_1228 : _GEN_819; // @[LoadStoreQueue.scala 150:36]
  wire [1:0] _GEN_1346 = EntryValid_1 ? _GEN_1229 : _GEN_820; // @[LoadStoreQueue.scala 150:36]
  wire [1:0] _GEN_1347 = EntryValid_1 ? _GEN_1230 : _GEN_821; // @[LoadStoreQueue.scala 150:36]
  wire [1:0] _GEN_1348 = EntryValid_1 ? _GEN_1231 : _GEN_822; // @[LoadStoreQueue.scala 150:36]
  wire [1:0] _GEN_1349 = EntryValid_1 ? _GEN_1232 : _GEN_823; // @[LoadStoreQueue.scala 150:36]
  wire [1:0] _GEN_1350 = EntryValid_1 ? _GEN_1233 : _GEN_824; // @[LoadStoreQueue.scala 150:36]
  wire [1:0] _GEN_1351 = EntryValid_1 ? _GEN_1234 : _GEN_825; // @[LoadStoreQueue.scala 150:36]
  wire [1:0] _GEN_1352 = EntryValid_1 ? _GEN_1235 : _GEN_826; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1353 = EntryValid_1 ? _GEN_1236 : _GEN_827; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1354 = EntryValid_1 ? _GEN_1237 : _GEN_828; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1355 = EntryValid_1 ? _GEN_1238 : _GEN_829; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1356 = EntryValid_1 ? _GEN_1239 : _GEN_830; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1357 = EntryValid_1 ? _GEN_1240 : _GEN_831; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1358 = EntryValid_1 ? _GEN_1241 : _GEN_832; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1359 = EntryValid_1 ? _GEN_1242 : _GEN_833; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1360 = EntryValid_1 ? _GEN_1243 : _GEN_834; // @[LoadStoreQueue.scala 150:36]
  wire [3:0] _GEN_1361 = EntryValid_1 ? _GEN_1244 : _GEN_835; // @[LoadStoreQueue.scala 150:36]
  wire [3:0] _GEN_1362 = EntryValid_1 ? _GEN_1245 : _GEN_836; // @[LoadStoreQueue.scala 150:36]
  wire [3:0] _GEN_1363 = EntryValid_1 ? _GEN_1246 : _GEN_837; // @[LoadStoreQueue.scala 150:36]
  wire [3:0] _GEN_1364 = EntryValid_1 ? _GEN_1247 : _GEN_838; // @[LoadStoreQueue.scala 150:36]
  wire [3:0] _GEN_1365 = EntryValid_1 ? _GEN_1248 : _GEN_839; // @[LoadStoreQueue.scala 150:36]
  wire [3:0] _GEN_1366 = EntryValid_1 ? _GEN_1249 : _GEN_840; // @[LoadStoreQueue.scala 150:36]
  wire [3:0] _GEN_1367 = EntryValid_1 ? _GEN_1250 : _GEN_841; // @[LoadStoreQueue.scala 150:36]
  wire [3:0] _GEN_1368 = EntryValid_1 ? _GEN_1251 : _GEN_842; // @[LoadStoreQueue.scala 150:36]
  wire [63:0] _GEN_1369 = EntryValid_1 ? _GEN_1252 : _GEN_843; // @[LoadStoreQueue.scala 150:36]
  wire [63:0] _GEN_1370 = EntryValid_1 ? _GEN_1253 : _GEN_844; // @[LoadStoreQueue.scala 150:36]
  wire [63:0] _GEN_1371 = EntryValid_1 ? _GEN_1254 : _GEN_845; // @[LoadStoreQueue.scala 150:36]
  wire [63:0] _GEN_1372 = EntryValid_1 ? _GEN_1255 : _GEN_846; // @[LoadStoreQueue.scala 150:36]
  wire [63:0] _GEN_1373 = EntryValid_1 ? _GEN_1256 : _GEN_847; // @[LoadStoreQueue.scala 150:36]
  wire [63:0] _GEN_1374 = EntryValid_1 ? _GEN_1257 : _GEN_848; // @[LoadStoreQueue.scala 150:36]
  wire [63:0] _GEN_1375 = EntryValid_1 ? _GEN_1258 : _GEN_849; // @[LoadStoreQueue.scala 150:36]
  wire [63:0] _GEN_1376 = EntryValid_1 ? _GEN_1259 : _GEN_850; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1377 = EntryValid_1 ? _GEN_1260 : _GEN_851; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1378 = EntryValid_1 ? _GEN_1261 : _GEN_852; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1379 = EntryValid_1 ? _GEN_1262 : _GEN_853; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1380 = EntryValid_1 ? _GEN_1263 : _GEN_854; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1381 = EntryValid_1 ? _GEN_1264 : _GEN_855; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1382 = EntryValid_1 ? _GEN_1265 : _GEN_856; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1383 = EntryValid_1 ? _GEN_1266 : _GEN_857; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1384 = EntryValid_1 ? _GEN_1267 : _GEN_858; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1385 = EntryValid_1 ? _GEN_1268 : _GEN_859; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1386 = EntryValid_1 ? _GEN_1269 : _GEN_860; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1387 = EntryValid_1 ? _GEN_1270 : _GEN_861; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1388 = EntryValid_1 ? _GEN_1271 : _GEN_862; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1389 = EntryValid_1 ? _GEN_1272 : _GEN_863; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1390 = EntryValid_1 ? _GEN_1273 : _GEN_864; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1391 = EntryValid_1 ? _GEN_1274 : _GEN_865; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1392 = EntryValid_1 ? _GEN_1275 : _GEN_866; // @[LoadStoreQueue.scala 150:36]
  wire [3:0] _GEN_1393 = EntryValid_1 ? _GEN_1276 : _GEN_867; // @[LoadStoreQueue.scala 150:36]
  wire [3:0] _GEN_1394 = EntryValid_1 ? _GEN_1277 : _GEN_868; // @[LoadStoreQueue.scala 150:36]
  wire [3:0] _GEN_1395 = EntryValid_1 ? _GEN_1278 : _GEN_869; // @[LoadStoreQueue.scala 150:36]
  wire [3:0] _GEN_1396 = EntryValid_1 ? _GEN_1279 : _GEN_870; // @[LoadStoreQueue.scala 150:36]
  wire [3:0] _GEN_1397 = EntryValid_1 ? _GEN_1280 : _GEN_871; // @[LoadStoreQueue.scala 150:36]
  wire [3:0] _GEN_1398 = EntryValid_1 ? _GEN_1281 : _GEN_872; // @[LoadStoreQueue.scala 150:36]
  wire [3:0] _GEN_1399 = EntryValid_1 ? _GEN_1282 : _GEN_873; // @[LoadStoreQueue.scala 150:36]
  wire [3:0] _GEN_1400 = EntryValid_1 ? _GEN_1283 : _GEN_874; // @[LoadStoreQueue.scala 150:36]
  wire [63:0] _GEN_1401 = EntryValid_1 ? _GEN_1284 : _GEN_875; // @[LoadStoreQueue.scala 150:36]
  wire [63:0] _GEN_1402 = EntryValid_1 ? _GEN_1285 : _GEN_876; // @[LoadStoreQueue.scala 150:36]
  wire [63:0] _GEN_1403 = EntryValid_1 ? _GEN_1286 : _GEN_877; // @[LoadStoreQueue.scala 150:36]
  wire [63:0] _GEN_1404 = EntryValid_1 ? _GEN_1287 : _GEN_878; // @[LoadStoreQueue.scala 150:36]
  wire [63:0] _GEN_1405 = EntryValid_1 ? _GEN_1288 : _GEN_879; // @[LoadStoreQueue.scala 150:36]
  wire [63:0] _GEN_1406 = EntryValid_1 ? _GEN_1289 : _GEN_880; // @[LoadStoreQueue.scala 150:36]
  wire [63:0] _GEN_1407 = EntryValid_1 ? _GEN_1290 : _GEN_881; // @[LoadStoreQueue.scala 150:36]
  wire [63:0] _GEN_1408 = EntryValid_1 ? _GEN_1291 : _GEN_882; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1409 = EntryValid_1 ? _GEN_1292 : _GEN_883; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1410 = EntryValid_1 ? _GEN_1293 : _GEN_884; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1411 = EntryValid_1 ? _GEN_1294 : _GEN_885; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1412 = EntryValid_1 ? _GEN_1295 : _GEN_886; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1413 = EntryValid_1 ? _GEN_1296 : _GEN_887; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1414 = EntryValid_1 ? _GEN_1297 : _GEN_888; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1415 = EntryValid_1 ? _GEN_1298 : _GEN_889; // @[LoadStoreQueue.scala 150:36]
  wire  _GEN_1416 = EntryValid_1 ? _GEN_1299 : _GEN_890; // @[LoadStoreQueue.scala 150:36]
  wire  _T_242 = checkOk | checkOk_1; // @[LoadStoreQueue.scala 192:19]
  wire [2:0] checkIndex_2 = nextTail + 3'h2; // @[LoadStoreQueue.scala 148:27]
  wire  _GEN_1418 = 3'h1 == checkIndex_2 ? buffer_1_valid : buffer_0_valid; // @[LoadStoreQueue.scala 150:{36,36}]
  wire  _GEN_1419 = 3'h2 == checkIndex_2 ? buffer_2_valid : _GEN_1418; // @[LoadStoreQueue.scala 150:{36,36}]
  wire  _GEN_1420 = 3'h3 == checkIndex_2 ? buffer_3_valid : _GEN_1419; // @[LoadStoreQueue.scala 150:{36,36}]
  wire  _GEN_1421 = 3'h4 == checkIndex_2 ? buffer_4_valid : _GEN_1420; // @[LoadStoreQueue.scala 150:{36,36}]
  wire  _GEN_1422 = 3'h5 == checkIndex_2 ? buffer_5_valid : _GEN_1421; // @[LoadStoreQueue.scala 150:{36,36}]
  wire  _GEN_1423 = 3'h6 == checkIndex_2 ? buffer_6_valid : _GEN_1422; // @[LoadStoreQueue.scala 150:{36,36}]
  wire  EntryValid_2 = 3'h7 == checkIndex_2 ? buffer_7_valid : _GEN_1423; // @[LoadStoreQueue.scala 150:{36,36}]
  wire [63:0] _GEN_1426 = 3'h1 == checkIndex_2 ? buffer_1_address : buffer_0_address; // @[LoadStoreQueue.scala 151:{18,18}]
  wire [63:0] _GEN_1427 = 3'h2 == checkIndex_2 ? buffer_2_address : _GEN_1426; // @[LoadStoreQueue.scala 151:{18,18}]
  wire [63:0] _GEN_1428 = 3'h3 == checkIndex_2 ? buffer_3_address : _GEN_1427; // @[LoadStoreQueue.scala 151:{18,18}]
  wire [63:0] _GEN_1429 = 3'h4 == checkIndex_2 ? buffer_4_address : _GEN_1428; // @[LoadStoreQueue.scala 151:{18,18}]
  wire [63:0] _GEN_1430 = 3'h5 == checkIndex_2 ? buffer_5_address : _GEN_1429; // @[LoadStoreQueue.scala 151:{18,18}]
  wire [63:0] _GEN_1431 = 3'h6 == checkIndex_2 ? buffer_6_address : _GEN_1430; // @[LoadStoreQueue.scala 151:{18,18}]
  wire [63:0] _GEN_1432 = 3'h7 == checkIndex_2 ? buffer_7_address : _GEN_1431; // @[LoadStoreQueue.scala 151:{18,18}]
  wire  _GEN_1434 = 3'h1 == checkIndex_2 ? buffer_1_addressValid : buffer_0_addressValid; // @[LoadStoreQueue.scala 152:{23,23}]
  wire  _GEN_1435 = 3'h2 == checkIndex_2 ? buffer_2_addressValid : _GEN_1434; // @[LoadStoreQueue.scala 152:{23,23}]
  wire  _GEN_1436 = 3'h3 == checkIndex_2 ? buffer_3_addressValid : _GEN_1435; // @[LoadStoreQueue.scala 152:{23,23}]
  wire  _GEN_1437 = 3'h4 == checkIndex_2 ? buffer_4_addressValid : _GEN_1436; // @[LoadStoreQueue.scala 152:{23,23}]
  wire  _GEN_1438 = 3'h5 == checkIndex_2 ? buffer_5_addressValid : _GEN_1437; // @[LoadStoreQueue.scala 152:{23,23}]
  wire  _GEN_1439 = 3'h6 == checkIndex_2 ? buffer_6_addressValid : _GEN_1438; // @[LoadStoreQueue.scala 152:{23,23}]
  wire  _GEN_1440 = 3'h7 == checkIndex_2 ? buffer_7_addressValid : _GEN_1439; // @[LoadStoreQueue.scala 152:{23,23}]
  wire  _T_244 = AddressValid_0 & Address_0 == _GEN_1432; // @[LoadStoreQueue.scala 160:32]
  wire  _T_246 = _T_244 | ~AddressValid_0; // @[LoadStoreQueue.scala 162:26]
  wire  _GEN_1442 = EntryValid_0 & _T_246; // @[LoadStoreQueue.scala 127:25 158:31]
  wire  _T_248 = AddressValid_1 & Address_1 == _GEN_1432; // @[LoadStoreQueue.scala 160:32]
  wire  _T_250 = _T_248 | ~AddressValid_1; // @[LoadStoreQueue.scala 162:26]
  wire  _GEN_1443 = _T_250 | _GEN_1442; // @[LoadStoreQueue.scala 163:15 164:26]
  wire  _GEN_1444 = EntryValid_1 ? _GEN_1443 : _GEN_1442; // @[LoadStoreQueue.scala 158:31]
  wire  _checkOk_T_24 = head != nextTail & EntryValid_2 & _GEN_1440; // @[LoadStoreQueue.scala 171:62]
  wire  _GEN_1446 = 3'h1 == checkIndex_2 ? buffer_1_info_accessType : buffer_0_info_accessType; // @[LoadStoreQueue.scala 174:{46,46}]
  wire  _GEN_1447 = 3'h2 == checkIndex_2 ? buffer_2_info_accessType : _GEN_1446; // @[LoadStoreQueue.scala 174:{46,46}]
  wire  _GEN_1448 = 3'h3 == checkIndex_2 ? buffer_3_info_accessType : _GEN_1447; // @[LoadStoreQueue.scala 174:{46,46}]
  wire  _GEN_1449 = 3'h4 == checkIndex_2 ? buffer_4_info_accessType : _GEN_1448; // @[LoadStoreQueue.scala 174:{46,46}]
  wire  _GEN_1450 = 3'h5 == checkIndex_2 ? buffer_5_info_accessType : _GEN_1449; // @[LoadStoreQueue.scala 174:{46,46}]
  wire  _GEN_1451 = 3'h6 == checkIndex_2 ? buffer_6_info_accessType : _GEN_1450; // @[LoadStoreQueue.scala 174:{46,46}]
  wire  _GEN_1452 = 3'h7 == checkIndex_2 ? buffer_7_info_accessType : _GEN_1451; // @[LoadStoreQueue.scala 174:{46,46}]
  wire  Overlap_2 = EntryValid_2 & _GEN_1444; // @[LoadStoreQueue.scala 127:25 150:36]
  wire  _GEN_1454 = 3'h1 == checkIndex_2 ? buffer_1_storeDataValid : buffer_0_storeDataValid; // @[LoadStoreQueue.scala 175:{57,57}]
  wire  _GEN_1455 = 3'h2 == checkIndex_2 ? buffer_2_storeDataValid : _GEN_1454; // @[LoadStoreQueue.scala 175:{57,57}]
  wire  _GEN_1456 = 3'h3 == checkIndex_2 ? buffer_3_storeDataValid : _GEN_1455; // @[LoadStoreQueue.scala 175:{57,57}]
  wire  _GEN_1457 = 3'h4 == checkIndex_2 ? buffer_4_storeDataValid : _GEN_1456; // @[LoadStoreQueue.scala 175:{57,57}]
  wire  _GEN_1458 = 3'h5 == checkIndex_2 ? buffer_5_storeDataValid : _GEN_1457; // @[LoadStoreQueue.scala 175:{57,57}]
  wire  _GEN_1459 = 3'h6 == checkIndex_2 ? buffer_6_storeDataValid : _GEN_1458; // @[LoadStoreQueue.scala 175:{57,57}]
  wire  _GEN_1460 = 3'h7 == checkIndex_2 ? buffer_7_storeDataValid : _GEN_1459; // @[LoadStoreQueue.scala 175:{57,57}]
  wire  _checkOk_T_29 = ~_GEN_1452 & _GEN_1460; // @[LoadStoreQueue.scala 175:57]
  wire  _GEN_1462 = 3'h1 == checkIndex_2 ? buffer_1_readyReorderSign : buffer_0_readyReorderSign; // @[LoadStoreQueue.scala 177:{28,28}]
  wire  _GEN_1463 = 3'h2 == checkIndex_2 ? buffer_2_readyReorderSign : _GEN_1462; // @[LoadStoreQueue.scala 177:{28,28}]
  wire  _GEN_1464 = 3'h3 == checkIndex_2 ? buffer_3_readyReorderSign : _GEN_1463; // @[LoadStoreQueue.scala 177:{28,28}]
  wire  _GEN_1465 = 3'h4 == checkIndex_2 ? buffer_4_readyReorderSign : _GEN_1464; // @[LoadStoreQueue.scala 177:{28,28}]
  wire  _GEN_1466 = 3'h5 == checkIndex_2 ? buffer_5_readyReorderSign : _GEN_1465; // @[LoadStoreQueue.scala 177:{28,28}]
  wire  _GEN_1467 = 3'h6 == checkIndex_2 ? buffer_6_readyReorderSign : _GEN_1466; // @[LoadStoreQueue.scala 177:{28,28}]
  wire  _GEN_1468 = 3'h7 == checkIndex_2 ? buffer_7_readyReorderSign : _GEN_1467; // @[LoadStoreQueue.scala 177:{28,28}]
  wire  _checkOk_T_30 = _checkOk_T_29 & _GEN_1468; // @[LoadStoreQueue.scala 177:28]
  wire  _checkOk_T_31 = _GEN_1452 & ~Overlap_2 | _checkOk_T_30; // @[LoadStoreQueue.scala 174:71]
  wire  _checkOk_T_32 = _checkOk_T_24 & _checkOk_T_31; // @[LoadStoreQueue.scala 173:22]
  wire  checkOk_2 = EntryValid_2 & _checkOk_T_32; // @[LoadStoreQueue.scala 150:36 171:15 149:30]
  wire  _GEN_1470 = 3'h1 == checkIndex_2 ? buffer_1_addressAndLoadResultTag_threadId :
    buffer_0_addressAndLoadResultTag_threadId; // @[LoadStoreQueue.scala 182:{28,28}]
  wire  _GEN_1471 = 3'h2 == checkIndex_2 ? buffer_2_addressAndLoadResultTag_threadId : _GEN_1470; // @[LoadStoreQueue.scala 182:{28,28}]
  wire  _GEN_1472 = 3'h3 == checkIndex_2 ? buffer_3_addressAndLoadResultTag_threadId : _GEN_1471; // @[LoadStoreQueue.scala 182:{28,28}]
  wire  _GEN_1473 = 3'h4 == checkIndex_2 ? buffer_4_addressAndLoadResultTag_threadId : _GEN_1472; // @[LoadStoreQueue.scala 182:{28,28}]
  wire  _GEN_1474 = 3'h5 == checkIndex_2 ? buffer_5_addressAndLoadResultTag_threadId : _GEN_1473; // @[LoadStoreQueue.scala 182:{28,28}]
  wire  _GEN_1475 = 3'h6 == checkIndex_2 ? buffer_6_addressAndLoadResultTag_threadId : _GEN_1474; // @[LoadStoreQueue.scala 182:{28,28}]
  wire  _GEN_1476 = 3'h7 == checkIndex_2 ? buffer_7_addressAndLoadResultTag_threadId : _GEN_1475; // @[LoadStoreQueue.scala 182:{28,28}]
  wire [3:0] _GEN_1478 = 3'h1 == checkIndex_2 ? buffer_1_addressAndLoadResultTag_id :
    buffer_0_addressAndLoadResultTag_id; // @[LoadStoreQueue.scala 182:{28,28}]
  wire [3:0] _GEN_1479 = 3'h2 == checkIndex_2 ? buffer_2_addressAndLoadResultTag_id : _GEN_1478; // @[LoadStoreQueue.scala 182:{28,28}]
  wire [3:0] _GEN_1480 = 3'h3 == checkIndex_2 ? buffer_3_addressAndLoadResultTag_id : _GEN_1479; // @[LoadStoreQueue.scala 182:{28,28}]
  wire [3:0] _GEN_1481 = 3'h4 == checkIndex_2 ? buffer_4_addressAndLoadResultTag_id : _GEN_1480; // @[LoadStoreQueue.scala 182:{28,28}]
  wire [3:0] _GEN_1482 = 3'h5 == checkIndex_2 ? buffer_5_addressAndLoadResultTag_id : _GEN_1481; // @[LoadStoreQueue.scala 182:{28,28}]
  wire [3:0] _GEN_1483 = 3'h6 == checkIndex_2 ? buffer_6_addressAndLoadResultTag_id : _GEN_1482; // @[LoadStoreQueue.scala 182:{28,28}]
  wire [3:0] _GEN_1484 = 3'h7 == checkIndex_2 ? buffer_7_addressAndLoadResultTag_id : _GEN_1483; // @[LoadStoreQueue.scala 182:{28,28}]
  wire [63:0] _GEN_1486 = 3'h1 == checkIndex_2 ? buffer_1_storeData : buffer_0_storeData; // @[LoadStoreQueue.scala 183:{29,29}]
  wire [63:0] _GEN_1487 = 3'h2 == checkIndex_2 ? buffer_2_storeData : _GEN_1486; // @[LoadStoreQueue.scala 183:{29,29}]
  wire [63:0] _GEN_1488 = 3'h3 == checkIndex_2 ? buffer_3_storeData : _GEN_1487; // @[LoadStoreQueue.scala 183:{29,29}]
  wire [63:0] _GEN_1489 = 3'h4 == checkIndex_2 ? buffer_4_storeData : _GEN_1488; // @[LoadStoreQueue.scala 183:{29,29}]
  wire [63:0] _GEN_1490 = 3'h5 == checkIndex_2 ? buffer_5_storeData : _GEN_1489; // @[LoadStoreQueue.scala 183:{29,29}]
  wire [63:0] _GEN_1491 = 3'h6 == checkIndex_2 ? buffer_6_storeData : _GEN_1490; // @[LoadStoreQueue.scala 183:{29,29}]
  wire [63:0] _GEN_1492 = 3'h7 == checkIndex_2 ? buffer_7_storeData : _GEN_1491; // @[LoadStoreQueue.scala 183:{29,29}]
  wire  _GEN_1494 = 3'h1 == checkIndex_2 ? buffer_1_info_signed : buffer_0_info_signed; // @[LoadStoreQueue.scala 185:{35,35}]
  wire  _GEN_1495 = 3'h2 == checkIndex_2 ? buffer_2_info_signed : _GEN_1494; // @[LoadStoreQueue.scala 185:{35,35}]
  wire  _GEN_1496 = 3'h3 == checkIndex_2 ? buffer_3_info_signed : _GEN_1495; // @[LoadStoreQueue.scala 185:{35,35}]
  wire  _GEN_1497 = 3'h4 == checkIndex_2 ? buffer_4_info_signed : _GEN_1496; // @[LoadStoreQueue.scala 185:{35,35}]
  wire  _GEN_1498 = 3'h5 == checkIndex_2 ? buffer_5_info_signed : _GEN_1497; // @[LoadStoreQueue.scala 185:{35,35}]
  wire  _GEN_1499 = 3'h6 == checkIndex_2 ? buffer_6_info_signed : _GEN_1498; // @[LoadStoreQueue.scala 185:{35,35}]
  wire  _GEN_1500 = 3'h7 == checkIndex_2 ? buffer_7_info_signed : _GEN_1499; // @[LoadStoreQueue.scala 185:{35,35}]
  wire [1:0] _GEN_1502 = 3'h1 == checkIndex_2 ? buffer_1_info_accessWidth : buffer_0_info_accessWidth; // @[LoadStoreQueue.scala 185:{35,35}]
  wire [1:0] _GEN_1503 = 3'h2 == checkIndex_2 ? buffer_2_info_accessWidth : _GEN_1502; // @[LoadStoreQueue.scala 185:{35,35}]
  wire [1:0] _GEN_1504 = 3'h3 == checkIndex_2 ? buffer_3_info_accessWidth : _GEN_1503; // @[LoadStoreQueue.scala 185:{35,35}]
  wire [1:0] _GEN_1505 = 3'h4 == checkIndex_2 ? buffer_4_info_accessWidth : _GEN_1504; // @[LoadStoreQueue.scala 185:{35,35}]
  wire [1:0] _GEN_1506 = 3'h5 == checkIndex_2 ? buffer_5_info_accessWidth : _GEN_1505; // @[LoadStoreQueue.scala 185:{35,35}]
  wire [1:0] _GEN_1507 = 3'h6 == checkIndex_2 ? buffer_6_info_accessWidth : _GEN_1506; // @[LoadStoreQueue.scala 185:{35,35}]
  wire [1:0] _GEN_1508 = 3'h7 == checkIndex_2 ? buffer_7_info_accessWidth : _GEN_1507; // @[LoadStoreQueue.scala 185:{35,35}]
  wire  _GEN_1509 = 3'h0 == checkIndex_2 ? 1'h0 : _GEN_1313; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1510 = 3'h1 == checkIndex_2 ? 1'h0 : _GEN_1314; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1511 = 3'h2 == checkIndex_2 ? 1'h0 : _GEN_1315; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1512 = 3'h3 == checkIndex_2 ? 1'h0 : _GEN_1316; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1513 = 3'h4 == checkIndex_2 ? 1'h0 : _GEN_1317; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1514 = 3'h5 == checkIndex_2 ? 1'h0 : _GEN_1318; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1515 = 3'h6 == checkIndex_2 ? 1'h0 : _GEN_1319; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1516 = 3'h7 == checkIndex_2 ? 1'h0 : _GEN_1320; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1517 = 3'h0 == checkIndex_2 ? 1'h0 : _GEN_1321; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1518 = 3'h1 == checkIndex_2 ? 1'h0 : _GEN_1322; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1519 = 3'h2 == checkIndex_2 ? 1'h0 : _GEN_1323; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1520 = 3'h3 == checkIndex_2 ? 1'h0 : _GEN_1324; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1521 = 3'h4 == checkIndex_2 ? 1'h0 : _GEN_1325; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1522 = 3'h5 == checkIndex_2 ? 1'h0 : _GEN_1326; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1523 = 3'h6 == checkIndex_2 ? 1'h0 : _GEN_1327; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1524 = 3'h7 == checkIndex_2 ? 1'h0 : _GEN_1328; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1549 = 3'h0 == checkIndex_2 ? 1'h0 : _GEN_1353; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1550 = 3'h1 == checkIndex_2 ? 1'h0 : _GEN_1354; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1551 = 3'h2 == checkIndex_2 ? 1'h0 : _GEN_1355; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1552 = 3'h3 == checkIndex_2 ? 1'h0 : _GEN_1356; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1553 = 3'h4 == checkIndex_2 ? 1'h0 : _GEN_1357; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1554 = 3'h5 == checkIndex_2 ? 1'h0 : _GEN_1358; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1555 = 3'h6 == checkIndex_2 ? 1'h0 : _GEN_1359; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1556 = 3'h7 == checkIndex_2 ? 1'h0 : _GEN_1360; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [3:0] _GEN_1557 = 3'h0 == checkIndex_2 ? 4'h0 : _GEN_1361; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [3:0] _GEN_1558 = 3'h1 == checkIndex_2 ? 4'h0 : _GEN_1362; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [3:0] _GEN_1559 = 3'h2 == checkIndex_2 ? 4'h0 : _GEN_1363; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [3:0] _GEN_1560 = 3'h3 == checkIndex_2 ? 4'h0 : _GEN_1364; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [3:0] _GEN_1561 = 3'h4 == checkIndex_2 ? 4'h0 : _GEN_1365; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [3:0] _GEN_1562 = 3'h5 == checkIndex_2 ? 4'h0 : _GEN_1366; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [3:0] _GEN_1563 = 3'h6 == checkIndex_2 ? 4'h0 : _GEN_1367; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [3:0] _GEN_1564 = 3'h7 == checkIndex_2 ? 4'h0 : _GEN_1368; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [63:0] _GEN_1565 = 3'h0 == checkIndex_2 ? 64'h0 : _GEN_1369; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [63:0] _GEN_1566 = 3'h1 == checkIndex_2 ? 64'h0 : _GEN_1370; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [63:0] _GEN_1567 = 3'h2 == checkIndex_2 ? 64'h0 : _GEN_1371; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [63:0] _GEN_1568 = 3'h3 == checkIndex_2 ? 64'h0 : _GEN_1372; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [63:0] _GEN_1569 = 3'h4 == checkIndex_2 ? 64'h0 : _GEN_1373; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [63:0] _GEN_1570 = 3'h5 == checkIndex_2 ? 64'h0 : _GEN_1374; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [63:0] _GEN_1571 = 3'h6 == checkIndex_2 ? 64'h0 : _GEN_1375; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [63:0] _GEN_1572 = 3'h7 == checkIndex_2 ? 64'h0 : _GEN_1376; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1573 = 3'h0 == checkIndex_2 ? 1'h0 : _GEN_1377; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1574 = 3'h1 == checkIndex_2 ? 1'h0 : _GEN_1378; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1575 = 3'h2 == checkIndex_2 ? 1'h0 : _GEN_1379; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1576 = 3'h3 == checkIndex_2 ? 1'h0 : _GEN_1380; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1577 = 3'h4 == checkIndex_2 ? 1'h0 : _GEN_1381; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1578 = 3'h5 == checkIndex_2 ? 1'h0 : _GEN_1382; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1579 = 3'h6 == checkIndex_2 ? 1'h0 : _GEN_1383; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1580 = 3'h7 == checkIndex_2 ? 1'h0 : _GEN_1384; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1581 = 3'h0 == checkIndex_2 ? 1'h0 : _GEN_1385; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1582 = 3'h1 == checkIndex_2 ? 1'h0 : _GEN_1386; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1583 = 3'h2 == checkIndex_2 ? 1'h0 : _GEN_1387; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1584 = 3'h3 == checkIndex_2 ? 1'h0 : _GEN_1388; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1585 = 3'h4 == checkIndex_2 ? 1'h0 : _GEN_1389; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1586 = 3'h5 == checkIndex_2 ? 1'h0 : _GEN_1390; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1587 = 3'h6 == checkIndex_2 ? 1'h0 : _GEN_1391; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1588 = 3'h7 == checkIndex_2 ? 1'h0 : _GEN_1392; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [3:0] _GEN_1589 = 3'h0 == checkIndex_2 ? 4'h0 : _GEN_1393; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [3:0] _GEN_1590 = 3'h1 == checkIndex_2 ? 4'h0 : _GEN_1394; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [3:0] _GEN_1591 = 3'h2 == checkIndex_2 ? 4'h0 : _GEN_1395; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [3:0] _GEN_1592 = 3'h3 == checkIndex_2 ? 4'h0 : _GEN_1396; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [3:0] _GEN_1593 = 3'h4 == checkIndex_2 ? 4'h0 : _GEN_1397; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [3:0] _GEN_1594 = 3'h5 == checkIndex_2 ? 4'h0 : _GEN_1398; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [3:0] _GEN_1595 = 3'h6 == checkIndex_2 ? 4'h0 : _GEN_1399; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [3:0] _GEN_1596 = 3'h7 == checkIndex_2 ? 4'h0 : _GEN_1400; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [63:0] _GEN_1597 = 3'h0 == checkIndex_2 ? 64'h0 : _GEN_1401; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [63:0] _GEN_1598 = 3'h1 == checkIndex_2 ? 64'h0 : _GEN_1402; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [63:0] _GEN_1599 = 3'h2 == checkIndex_2 ? 64'h0 : _GEN_1403; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [63:0] _GEN_1600 = 3'h3 == checkIndex_2 ? 64'h0 : _GEN_1404; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [63:0] _GEN_1601 = 3'h4 == checkIndex_2 ? 64'h0 : _GEN_1405; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [63:0] _GEN_1602 = 3'h5 == checkIndex_2 ? 64'h0 : _GEN_1406; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [63:0] _GEN_1603 = 3'h6 == checkIndex_2 ? 64'h0 : _GEN_1407; // @[LoadStoreQueue.scala 187:{30,30}]
  wire [63:0] _GEN_1604 = 3'h7 == checkIndex_2 ? 64'h0 : _GEN_1408; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1605 = 3'h0 == checkIndex_2 ? 1'h0 : _GEN_1409; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1606 = 3'h1 == checkIndex_2 ? 1'h0 : _GEN_1410; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1607 = 3'h2 == checkIndex_2 ? 1'h0 : _GEN_1411; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1608 = 3'h3 == checkIndex_2 ? 1'h0 : _GEN_1412; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1609 = 3'h4 == checkIndex_2 ? 1'h0 : _GEN_1413; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1610 = 3'h5 == checkIndex_2 ? 1'h0 : _GEN_1414; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1611 = 3'h6 == checkIndex_2 ? 1'h0 : _GEN_1415; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1612 = 3'h7 == checkIndex_2 ? 1'h0 : _GEN_1416; // @[LoadStoreQueue.scala 187:{30,30}]
  wire  _GEN_1717 = checkOk_2 & ~_T_242 ? _GEN_1476 : _GEN_1306; // @[LoadStoreQueue.scala 181:31 182:28]
  wire [3:0] _GEN_1718 = checkOk_2 & ~_T_242 ? _GEN_1484 : _GEN_1307; // @[LoadStoreQueue.scala 181:31 182:28]
  wire [63:0] _GEN_1719 = checkOk_2 & ~_T_242 ? _GEN_1492 : _GEN_1308; // @[LoadStoreQueue.scala 181:31 183:29]
  wire [63:0] _GEN_1720 = checkOk_2 & ~_T_242 ? _GEN_1432 : _GEN_1309; // @[LoadStoreQueue.scala 181:31 184:32]
  wire  _GEN_1721 = checkOk_2 & ~_T_242 ? _GEN_1452 : _GEN_1310; // @[LoadStoreQueue.scala 181:31 185:35]
  wire  _GEN_1722 = checkOk_2 & ~_T_242 ? _GEN_1500 : _GEN_1311; // @[LoadStoreQueue.scala 181:31 185:35]
  wire [1:0] _GEN_1723 = checkOk_2 & ~_T_242 ? _GEN_1508 : _GEN_1312; // @[LoadStoreQueue.scala 181:31 185:35]
  wire  _GEN_1946 = 3'h1 == nextTail ? buffer_1_valid : buffer_0_valid; // @[LoadStoreQueue.scala 194:{8,8}]
  wire  _GEN_1947 = 3'h2 == nextTail ? buffer_2_valid : _GEN_1946; // @[LoadStoreQueue.scala 194:{8,8}]
  wire  _GEN_1948 = 3'h3 == nextTail ? buffer_3_valid : _GEN_1947; // @[LoadStoreQueue.scala 194:{8,8}]
  wire  _GEN_1949 = 3'h4 == nextTail ? buffer_4_valid : _GEN_1948; // @[LoadStoreQueue.scala 194:{8,8}]
  wire  _GEN_1950 = 3'h5 == nextTail ? buffer_5_valid : _GEN_1949; // @[LoadStoreQueue.scala 194:{8,8}]
  wire  _GEN_1951 = 3'h6 == nextTail ? buffer_6_valid : _GEN_1950; // @[LoadStoreQueue.scala 194:{8,8}]
  wire  _GEN_1952 = 3'h7 == nextTail ? buffer_7_valid : _GEN_1951; // @[LoadStoreQueue.scala 194:{8,8}]
  assign io_decoders_0_ready = nextTail != _io_decoders_0_ready_T_1; // @[LoadStoreQueue.scala 61:27]
  assign io_memory_valid = EntryValid_2 ? checkOk_2 | _T_242 : _GEN_1305; // @[LoadStoreQueue.scala 150:36 179:23]
  assign io_memory_bits_address = EntryValid_2 ? _GEN_1720 : _GEN_1309; // @[LoadStoreQueue.scala 150:36]
  assign io_memory_bits_tag_threadId = EntryValid_2 ? _GEN_1717 : _GEN_1306; // @[LoadStoreQueue.scala 150:36]
  assign io_memory_bits_tag_id = EntryValid_2 ? _GEN_1718 : _GEN_1307; // @[LoadStoreQueue.scala 150:36]
  assign io_memory_bits_data = EntryValid_2 ? _GEN_1719 : _GEN_1308; // @[LoadStoreQueue.scala 150:36]
  assign io_memory_bits_accessInfo_accessType = EntryValid_2 ? _GEN_1721 : _GEN_1310; // @[LoadStoreQueue.scala 150:36]
  assign io_memory_bits_accessInfo_signed = EntryValid_2 ? _GEN_1722 : _GEN_1311; // @[LoadStoreQueue.scala 150:36]
  assign io_memory_bits_accessInfo_accessWidth = EntryValid_2 ? _GEN_1723 : _GEN_1312; // @[LoadStoreQueue.scala 150:36]
  assign io_isEmpty = head == nextTail; // @[LoadStoreQueue.scala 49:22]
  always @(posedge clock) begin
    if (reset) begin // @[LoadStoreQueue.scala 47:21]
      head <= 3'h0; // @[LoadStoreQueue.scala 47:21]
    end else begin
      head <= insertIndex; // @[LoadStoreQueue.scala 84:8]
    end
    if (reset) begin // @[LoadStoreQueue.scala 48:21]
      nextTail <= 3'h0; // @[LoadStoreQueue.scala 48:21]
    end else if (~_GEN_1952 & _checkOk_T) begin // @[LoadStoreQueue.scala 194:46]
      nextTail <= checkIndex_1; // @[LoadStoreQueue.scala 195:10]
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_0_valid <= 1'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_0_valid <= _GEN_1509;
        end else begin
          buffer_0_valid <= _GEN_1313;
        end
      end else begin
        buffer_0_valid <= _GEN_1313;
      end
    end else begin
      buffer_0_valid <= _GEN_1313;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_0_readyReorderSign <= 1'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_0_readyReorderSign <= _GEN_1517;
        end else begin
          buffer_0_readyReorderSign <= _GEN_1321;
        end
      end else begin
        buffer_0_readyReorderSign <= _GEN_1321;
      end
    end else begin
      buffer_0_readyReorderSign <= _GEN_1321;
    end
    if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          if (3'h0 == checkIndex_2) begin // @[LoadStoreQueue.scala 187:30]
            buffer_0_info_accessType <= 1'h0; // @[LoadStoreQueue.scala 187:30]
          end else begin
            buffer_0_info_accessType <= _GEN_1329;
          end
        end else begin
          buffer_0_info_accessType <= _GEN_1329;
        end
      end else begin
        buffer_0_info_accessType <= _GEN_1329;
      end
    end else begin
      buffer_0_info_accessType <= _GEN_1329;
    end
    if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          if (3'h0 == checkIndex_2) begin // @[LoadStoreQueue.scala 187:30]
            buffer_0_info_signed <= 1'h0; // @[LoadStoreQueue.scala 187:30]
          end else begin
            buffer_0_info_signed <= _GEN_1337;
          end
        end else begin
          buffer_0_info_signed <= _GEN_1337;
        end
      end else begin
        buffer_0_info_signed <= _GEN_1337;
      end
    end else begin
      buffer_0_info_signed <= _GEN_1337;
    end
    if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          if (3'h0 == checkIndex_2) begin // @[LoadStoreQueue.scala 187:30]
            buffer_0_info_accessWidth <= 2'h0; // @[LoadStoreQueue.scala 187:30]
          end else begin
            buffer_0_info_accessWidth <= _GEN_1345;
          end
        end else begin
          buffer_0_info_accessWidth <= _GEN_1345;
        end
      end else begin
        buffer_0_info_accessWidth <= _GEN_1345;
      end
    end else begin
      buffer_0_info_accessWidth <= _GEN_1345;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_0_addressAndLoadResultTag_threadId <= 1'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_0_addressAndLoadResultTag_threadId <= _GEN_1549;
        end else begin
          buffer_0_addressAndLoadResultTag_threadId <= _GEN_1353;
        end
      end else begin
        buffer_0_addressAndLoadResultTag_threadId <= _GEN_1353;
      end
    end else begin
      buffer_0_addressAndLoadResultTag_threadId <= _GEN_1353;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_0_addressAndLoadResultTag_id <= 4'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_0_addressAndLoadResultTag_id <= _GEN_1557;
        end else begin
          buffer_0_addressAndLoadResultTag_id <= _GEN_1361;
        end
      end else begin
        buffer_0_addressAndLoadResultTag_id <= _GEN_1361;
      end
    end else begin
      buffer_0_addressAndLoadResultTag_id <= _GEN_1361;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_0_address <= 64'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_0_address <= _GEN_1565;
        end else begin
          buffer_0_address <= _GEN_1369;
        end
      end else begin
        buffer_0_address <= _GEN_1369;
      end
    end else begin
      buffer_0_address <= _GEN_1369;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_0_addressValid <= 1'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_0_addressValid <= _GEN_1573;
        end else begin
          buffer_0_addressValid <= _GEN_1377;
        end
      end else begin
        buffer_0_addressValid <= _GEN_1377;
      end
    end else begin
      buffer_0_addressValid <= _GEN_1377;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_0_storeDataTag_threadId <= 1'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_0_storeDataTag_threadId <= _GEN_1581;
        end else begin
          buffer_0_storeDataTag_threadId <= _GEN_1385;
        end
      end else begin
        buffer_0_storeDataTag_threadId <= _GEN_1385;
      end
    end else begin
      buffer_0_storeDataTag_threadId <= _GEN_1385;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_0_storeDataTag_id <= 4'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_0_storeDataTag_id <= _GEN_1589;
        end else begin
          buffer_0_storeDataTag_id <= _GEN_1393;
        end
      end else begin
        buffer_0_storeDataTag_id <= _GEN_1393;
      end
    end else begin
      buffer_0_storeDataTag_id <= _GEN_1393;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_0_storeData <= 64'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_0_storeData <= _GEN_1597;
        end else begin
          buffer_0_storeData <= _GEN_1401;
        end
      end else begin
        buffer_0_storeData <= _GEN_1401;
      end
    end else begin
      buffer_0_storeData <= _GEN_1401;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_0_storeDataValid <= 1'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_0_storeDataValid <= _GEN_1605;
        end else begin
          buffer_0_storeDataValid <= _GEN_1409;
        end
      end else begin
        buffer_0_storeDataValid <= _GEN_1409;
      end
    end else begin
      buffer_0_storeDataValid <= _GEN_1409;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_1_valid <= 1'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_1_valid <= _GEN_1510;
        end else begin
          buffer_1_valid <= _GEN_1314;
        end
      end else begin
        buffer_1_valid <= _GEN_1314;
      end
    end else begin
      buffer_1_valid <= _GEN_1314;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_1_readyReorderSign <= 1'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_1_readyReorderSign <= _GEN_1518;
        end else begin
          buffer_1_readyReorderSign <= _GEN_1322;
        end
      end else begin
        buffer_1_readyReorderSign <= _GEN_1322;
      end
    end else begin
      buffer_1_readyReorderSign <= _GEN_1322;
    end
    if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          if (3'h1 == checkIndex_2) begin // @[LoadStoreQueue.scala 187:30]
            buffer_1_info_accessType <= 1'h0; // @[LoadStoreQueue.scala 187:30]
          end else begin
            buffer_1_info_accessType <= _GEN_1330;
          end
        end else begin
          buffer_1_info_accessType <= _GEN_1330;
        end
      end else begin
        buffer_1_info_accessType <= _GEN_1330;
      end
    end else begin
      buffer_1_info_accessType <= _GEN_1330;
    end
    if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          if (3'h1 == checkIndex_2) begin // @[LoadStoreQueue.scala 187:30]
            buffer_1_info_signed <= 1'h0; // @[LoadStoreQueue.scala 187:30]
          end else begin
            buffer_1_info_signed <= _GEN_1338;
          end
        end else begin
          buffer_1_info_signed <= _GEN_1338;
        end
      end else begin
        buffer_1_info_signed <= _GEN_1338;
      end
    end else begin
      buffer_1_info_signed <= _GEN_1338;
    end
    if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          if (3'h1 == checkIndex_2) begin // @[LoadStoreQueue.scala 187:30]
            buffer_1_info_accessWidth <= 2'h0; // @[LoadStoreQueue.scala 187:30]
          end else begin
            buffer_1_info_accessWidth <= _GEN_1346;
          end
        end else begin
          buffer_1_info_accessWidth <= _GEN_1346;
        end
      end else begin
        buffer_1_info_accessWidth <= _GEN_1346;
      end
    end else begin
      buffer_1_info_accessWidth <= _GEN_1346;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_1_addressAndLoadResultTag_threadId <= 1'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_1_addressAndLoadResultTag_threadId <= _GEN_1550;
        end else begin
          buffer_1_addressAndLoadResultTag_threadId <= _GEN_1354;
        end
      end else begin
        buffer_1_addressAndLoadResultTag_threadId <= _GEN_1354;
      end
    end else begin
      buffer_1_addressAndLoadResultTag_threadId <= _GEN_1354;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_1_addressAndLoadResultTag_id <= 4'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_1_addressAndLoadResultTag_id <= _GEN_1558;
        end else begin
          buffer_1_addressAndLoadResultTag_id <= _GEN_1362;
        end
      end else begin
        buffer_1_addressAndLoadResultTag_id <= _GEN_1362;
      end
    end else begin
      buffer_1_addressAndLoadResultTag_id <= _GEN_1362;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_1_address <= 64'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_1_address <= _GEN_1566;
        end else begin
          buffer_1_address <= _GEN_1370;
        end
      end else begin
        buffer_1_address <= _GEN_1370;
      end
    end else begin
      buffer_1_address <= _GEN_1370;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_1_addressValid <= 1'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_1_addressValid <= _GEN_1574;
        end else begin
          buffer_1_addressValid <= _GEN_1378;
        end
      end else begin
        buffer_1_addressValid <= _GEN_1378;
      end
    end else begin
      buffer_1_addressValid <= _GEN_1378;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_1_storeDataTag_threadId <= 1'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_1_storeDataTag_threadId <= _GEN_1582;
        end else begin
          buffer_1_storeDataTag_threadId <= _GEN_1386;
        end
      end else begin
        buffer_1_storeDataTag_threadId <= _GEN_1386;
      end
    end else begin
      buffer_1_storeDataTag_threadId <= _GEN_1386;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_1_storeDataTag_id <= 4'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_1_storeDataTag_id <= _GEN_1590;
        end else begin
          buffer_1_storeDataTag_id <= _GEN_1394;
        end
      end else begin
        buffer_1_storeDataTag_id <= _GEN_1394;
      end
    end else begin
      buffer_1_storeDataTag_id <= _GEN_1394;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_1_storeData <= 64'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_1_storeData <= _GEN_1598;
        end else begin
          buffer_1_storeData <= _GEN_1402;
        end
      end else begin
        buffer_1_storeData <= _GEN_1402;
      end
    end else begin
      buffer_1_storeData <= _GEN_1402;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_1_storeDataValid <= 1'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_1_storeDataValid <= _GEN_1606;
        end else begin
          buffer_1_storeDataValid <= _GEN_1410;
        end
      end else begin
        buffer_1_storeDataValid <= _GEN_1410;
      end
    end else begin
      buffer_1_storeDataValid <= _GEN_1410;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_2_valid <= 1'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_2_valid <= _GEN_1511;
        end else begin
          buffer_2_valid <= _GEN_1315;
        end
      end else begin
        buffer_2_valid <= _GEN_1315;
      end
    end else begin
      buffer_2_valid <= _GEN_1315;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_2_readyReorderSign <= 1'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_2_readyReorderSign <= _GEN_1519;
        end else begin
          buffer_2_readyReorderSign <= _GEN_1323;
        end
      end else begin
        buffer_2_readyReorderSign <= _GEN_1323;
      end
    end else begin
      buffer_2_readyReorderSign <= _GEN_1323;
    end
    if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          if (3'h2 == checkIndex_2) begin // @[LoadStoreQueue.scala 187:30]
            buffer_2_info_accessType <= 1'h0; // @[LoadStoreQueue.scala 187:30]
          end else begin
            buffer_2_info_accessType <= _GEN_1331;
          end
        end else begin
          buffer_2_info_accessType <= _GEN_1331;
        end
      end else begin
        buffer_2_info_accessType <= _GEN_1331;
      end
    end else begin
      buffer_2_info_accessType <= _GEN_1331;
    end
    if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          if (3'h2 == checkIndex_2) begin // @[LoadStoreQueue.scala 187:30]
            buffer_2_info_signed <= 1'h0; // @[LoadStoreQueue.scala 187:30]
          end else begin
            buffer_2_info_signed <= _GEN_1339;
          end
        end else begin
          buffer_2_info_signed <= _GEN_1339;
        end
      end else begin
        buffer_2_info_signed <= _GEN_1339;
      end
    end else begin
      buffer_2_info_signed <= _GEN_1339;
    end
    if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          if (3'h2 == checkIndex_2) begin // @[LoadStoreQueue.scala 187:30]
            buffer_2_info_accessWidth <= 2'h0; // @[LoadStoreQueue.scala 187:30]
          end else begin
            buffer_2_info_accessWidth <= _GEN_1347;
          end
        end else begin
          buffer_2_info_accessWidth <= _GEN_1347;
        end
      end else begin
        buffer_2_info_accessWidth <= _GEN_1347;
      end
    end else begin
      buffer_2_info_accessWidth <= _GEN_1347;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_2_addressAndLoadResultTag_threadId <= 1'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_2_addressAndLoadResultTag_threadId <= _GEN_1551;
        end else begin
          buffer_2_addressAndLoadResultTag_threadId <= _GEN_1355;
        end
      end else begin
        buffer_2_addressAndLoadResultTag_threadId <= _GEN_1355;
      end
    end else begin
      buffer_2_addressAndLoadResultTag_threadId <= _GEN_1355;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_2_addressAndLoadResultTag_id <= 4'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_2_addressAndLoadResultTag_id <= _GEN_1559;
        end else begin
          buffer_2_addressAndLoadResultTag_id <= _GEN_1363;
        end
      end else begin
        buffer_2_addressAndLoadResultTag_id <= _GEN_1363;
      end
    end else begin
      buffer_2_addressAndLoadResultTag_id <= _GEN_1363;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_2_address <= 64'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_2_address <= _GEN_1567;
        end else begin
          buffer_2_address <= _GEN_1371;
        end
      end else begin
        buffer_2_address <= _GEN_1371;
      end
    end else begin
      buffer_2_address <= _GEN_1371;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_2_addressValid <= 1'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_2_addressValid <= _GEN_1575;
        end else begin
          buffer_2_addressValid <= _GEN_1379;
        end
      end else begin
        buffer_2_addressValid <= _GEN_1379;
      end
    end else begin
      buffer_2_addressValid <= _GEN_1379;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_2_storeDataTag_threadId <= 1'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_2_storeDataTag_threadId <= _GEN_1583;
        end else begin
          buffer_2_storeDataTag_threadId <= _GEN_1387;
        end
      end else begin
        buffer_2_storeDataTag_threadId <= _GEN_1387;
      end
    end else begin
      buffer_2_storeDataTag_threadId <= _GEN_1387;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_2_storeDataTag_id <= 4'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_2_storeDataTag_id <= _GEN_1591;
        end else begin
          buffer_2_storeDataTag_id <= _GEN_1395;
        end
      end else begin
        buffer_2_storeDataTag_id <= _GEN_1395;
      end
    end else begin
      buffer_2_storeDataTag_id <= _GEN_1395;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_2_storeData <= 64'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_2_storeData <= _GEN_1599;
        end else begin
          buffer_2_storeData <= _GEN_1403;
        end
      end else begin
        buffer_2_storeData <= _GEN_1403;
      end
    end else begin
      buffer_2_storeData <= _GEN_1403;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_2_storeDataValid <= 1'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_2_storeDataValid <= _GEN_1607;
        end else begin
          buffer_2_storeDataValid <= _GEN_1411;
        end
      end else begin
        buffer_2_storeDataValid <= _GEN_1411;
      end
    end else begin
      buffer_2_storeDataValid <= _GEN_1411;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_3_valid <= 1'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_3_valid <= _GEN_1512;
        end else begin
          buffer_3_valid <= _GEN_1316;
        end
      end else begin
        buffer_3_valid <= _GEN_1316;
      end
    end else begin
      buffer_3_valid <= _GEN_1316;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_3_readyReorderSign <= 1'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_3_readyReorderSign <= _GEN_1520;
        end else begin
          buffer_3_readyReorderSign <= _GEN_1324;
        end
      end else begin
        buffer_3_readyReorderSign <= _GEN_1324;
      end
    end else begin
      buffer_3_readyReorderSign <= _GEN_1324;
    end
    if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          if (3'h3 == checkIndex_2) begin // @[LoadStoreQueue.scala 187:30]
            buffer_3_info_accessType <= 1'h0; // @[LoadStoreQueue.scala 187:30]
          end else begin
            buffer_3_info_accessType <= _GEN_1332;
          end
        end else begin
          buffer_3_info_accessType <= _GEN_1332;
        end
      end else begin
        buffer_3_info_accessType <= _GEN_1332;
      end
    end else begin
      buffer_3_info_accessType <= _GEN_1332;
    end
    if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          if (3'h3 == checkIndex_2) begin // @[LoadStoreQueue.scala 187:30]
            buffer_3_info_signed <= 1'h0; // @[LoadStoreQueue.scala 187:30]
          end else begin
            buffer_3_info_signed <= _GEN_1340;
          end
        end else begin
          buffer_3_info_signed <= _GEN_1340;
        end
      end else begin
        buffer_3_info_signed <= _GEN_1340;
      end
    end else begin
      buffer_3_info_signed <= _GEN_1340;
    end
    if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          if (3'h3 == checkIndex_2) begin // @[LoadStoreQueue.scala 187:30]
            buffer_3_info_accessWidth <= 2'h0; // @[LoadStoreQueue.scala 187:30]
          end else begin
            buffer_3_info_accessWidth <= _GEN_1348;
          end
        end else begin
          buffer_3_info_accessWidth <= _GEN_1348;
        end
      end else begin
        buffer_3_info_accessWidth <= _GEN_1348;
      end
    end else begin
      buffer_3_info_accessWidth <= _GEN_1348;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_3_addressAndLoadResultTag_threadId <= 1'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_3_addressAndLoadResultTag_threadId <= _GEN_1552;
        end else begin
          buffer_3_addressAndLoadResultTag_threadId <= _GEN_1356;
        end
      end else begin
        buffer_3_addressAndLoadResultTag_threadId <= _GEN_1356;
      end
    end else begin
      buffer_3_addressAndLoadResultTag_threadId <= _GEN_1356;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_3_addressAndLoadResultTag_id <= 4'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_3_addressAndLoadResultTag_id <= _GEN_1560;
        end else begin
          buffer_3_addressAndLoadResultTag_id <= _GEN_1364;
        end
      end else begin
        buffer_3_addressAndLoadResultTag_id <= _GEN_1364;
      end
    end else begin
      buffer_3_addressAndLoadResultTag_id <= _GEN_1364;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_3_address <= 64'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_3_address <= _GEN_1568;
        end else begin
          buffer_3_address <= _GEN_1372;
        end
      end else begin
        buffer_3_address <= _GEN_1372;
      end
    end else begin
      buffer_3_address <= _GEN_1372;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_3_addressValid <= 1'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_3_addressValid <= _GEN_1576;
        end else begin
          buffer_3_addressValid <= _GEN_1380;
        end
      end else begin
        buffer_3_addressValid <= _GEN_1380;
      end
    end else begin
      buffer_3_addressValid <= _GEN_1380;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_3_storeDataTag_threadId <= 1'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_3_storeDataTag_threadId <= _GEN_1584;
        end else begin
          buffer_3_storeDataTag_threadId <= _GEN_1388;
        end
      end else begin
        buffer_3_storeDataTag_threadId <= _GEN_1388;
      end
    end else begin
      buffer_3_storeDataTag_threadId <= _GEN_1388;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_3_storeDataTag_id <= 4'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_3_storeDataTag_id <= _GEN_1592;
        end else begin
          buffer_3_storeDataTag_id <= _GEN_1396;
        end
      end else begin
        buffer_3_storeDataTag_id <= _GEN_1396;
      end
    end else begin
      buffer_3_storeDataTag_id <= _GEN_1396;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_3_storeData <= 64'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_3_storeData <= _GEN_1600;
        end else begin
          buffer_3_storeData <= _GEN_1404;
        end
      end else begin
        buffer_3_storeData <= _GEN_1404;
      end
    end else begin
      buffer_3_storeData <= _GEN_1404;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_3_storeDataValid <= 1'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_3_storeDataValid <= _GEN_1608;
        end else begin
          buffer_3_storeDataValid <= _GEN_1412;
        end
      end else begin
        buffer_3_storeDataValid <= _GEN_1412;
      end
    end else begin
      buffer_3_storeDataValid <= _GEN_1412;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_4_valid <= 1'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_4_valid <= _GEN_1513;
        end else begin
          buffer_4_valid <= _GEN_1317;
        end
      end else begin
        buffer_4_valid <= _GEN_1317;
      end
    end else begin
      buffer_4_valid <= _GEN_1317;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_4_readyReorderSign <= 1'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_4_readyReorderSign <= _GEN_1521;
        end else begin
          buffer_4_readyReorderSign <= _GEN_1325;
        end
      end else begin
        buffer_4_readyReorderSign <= _GEN_1325;
      end
    end else begin
      buffer_4_readyReorderSign <= _GEN_1325;
    end
    if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          if (3'h4 == checkIndex_2) begin // @[LoadStoreQueue.scala 187:30]
            buffer_4_info_accessType <= 1'h0; // @[LoadStoreQueue.scala 187:30]
          end else begin
            buffer_4_info_accessType <= _GEN_1333;
          end
        end else begin
          buffer_4_info_accessType <= _GEN_1333;
        end
      end else begin
        buffer_4_info_accessType <= _GEN_1333;
      end
    end else begin
      buffer_4_info_accessType <= _GEN_1333;
    end
    if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          if (3'h4 == checkIndex_2) begin // @[LoadStoreQueue.scala 187:30]
            buffer_4_info_signed <= 1'h0; // @[LoadStoreQueue.scala 187:30]
          end else begin
            buffer_4_info_signed <= _GEN_1341;
          end
        end else begin
          buffer_4_info_signed <= _GEN_1341;
        end
      end else begin
        buffer_4_info_signed <= _GEN_1341;
      end
    end else begin
      buffer_4_info_signed <= _GEN_1341;
    end
    if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          if (3'h4 == checkIndex_2) begin // @[LoadStoreQueue.scala 187:30]
            buffer_4_info_accessWidth <= 2'h0; // @[LoadStoreQueue.scala 187:30]
          end else begin
            buffer_4_info_accessWidth <= _GEN_1349;
          end
        end else begin
          buffer_4_info_accessWidth <= _GEN_1349;
        end
      end else begin
        buffer_4_info_accessWidth <= _GEN_1349;
      end
    end else begin
      buffer_4_info_accessWidth <= _GEN_1349;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_4_addressAndLoadResultTag_threadId <= 1'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_4_addressAndLoadResultTag_threadId <= _GEN_1553;
        end else begin
          buffer_4_addressAndLoadResultTag_threadId <= _GEN_1357;
        end
      end else begin
        buffer_4_addressAndLoadResultTag_threadId <= _GEN_1357;
      end
    end else begin
      buffer_4_addressAndLoadResultTag_threadId <= _GEN_1357;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_4_addressAndLoadResultTag_id <= 4'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_4_addressAndLoadResultTag_id <= _GEN_1561;
        end else begin
          buffer_4_addressAndLoadResultTag_id <= _GEN_1365;
        end
      end else begin
        buffer_4_addressAndLoadResultTag_id <= _GEN_1365;
      end
    end else begin
      buffer_4_addressAndLoadResultTag_id <= _GEN_1365;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_4_address <= 64'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_4_address <= _GEN_1569;
        end else begin
          buffer_4_address <= _GEN_1373;
        end
      end else begin
        buffer_4_address <= _GEN_1373;
      end
    end else begin
      buffer_4_address <= _GEN_1373;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_4_addressValid <= 1'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_4_addressValid <= _GEN_1577;
        end else begin
          buffer_4_addressValid <= _GEN_1381;
        end
      end else begin
        buffer_4_addressValid <= _GEN_1381;
      end
    end else begin
      buffer_4_addressValid <= _GEN_1381;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_4_storeDataTag_threadId <= 1'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_4_storeDataTag_threadId <= _GEN_1585;
        end else begin
          buffer_4_storeDataTag_threadId <= _GEN_1389;
        end
      end else begin
        buffer_4_storeDataTag_threadId <= _GEN_1389;
      end
    end else begin
      buffer_4_storeDataTag_threadId <= _GEN_1389;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_4_storeDataTag_id <= 4'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_4_storeDataTag_id <= _GEN_1593;
        end else begin
          buffer_4_storeDataTag_id <= _GEN_1397;
        end
      end else begin
        buffer_4_storeDataTag_id <= _GEN_1397;
      end
    end else begin
      buffer_4_storeDataTag_id <= _GEN_1397;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_4_storeData <= 64'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_4_storeData <= _GEN_1601;
        end else begin
          buffer_4_storeData <= _GEN_1405;
        end
      end else begin
        buffer_4_storeData <= _GEN_1405;
      end
    end else begin
      buffer_4_storeData <= _GEN_1405;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_4_storeDataValid <= 1'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_4_storeDataValid <= _GEN_1609;
        end else begin
          buffer_4_storeDataValid <= _GEN_1413;
        end
      end else begin
        buffer_4_storeDataValid <= _GEN_1413;
      end
    end else begin
      buffer_4_storeDataValid <= _GEN_1413;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_5_valid <= 1'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_5_valid <= _GEN_1514;
        end else begin
          buffer_5_valid <= _GEN_1318;
        end
      end else begin
        buffer_5_valid <= _GEN_1318;
      end
    end else begin
      buffer_5_valid <= _GEN_1318;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_5_readyReorderSign <= 1'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_5_readyReorderSign <= _GEN_1522;
        end else begin
          buffer_5_readyReorderSign <= _GEN_1326;
        end
      end else begin
        buffer_5_readyReorderSign <= _GEN_1326;
      end
    end else begin
      buffer_5_readyReorderSign <= _GEN_1326;
    end
    if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          if (3'h5 == checkIndex_2) begin // @[LoadStoreQueue.scala 187:30]
            buffer_5_info_accessType <= 1'h0; // @[LoadStoreQueue.scala 187:30]
          end else begin
            buffer_5_info_accessType <= _GEN_1334;
          end
        end else begin
          buffer_5_info_accessType <= _GEN_1334;
        end
      end else begin
        buffer_5_info_accessType <= _GEN_1334;
      end
    end else begin
      buffer_5_info_accessType <= _GEN_1334;
    end
    if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          if (3'h5 == checkIndex_2) begin // @[LoadStoreQueue.scala 187:30]
            buffer_5_info_signed <= 1'h0; // @[LoadStoreQueue.scala 187:30]
          end else begin
            buffer_5_info_signed <= _GEN_1342;
          end
        end else begin
          buffer_5_info_signed <= _GEN_1342;
        end
      end else begin
        buffer_5_info_signed <= _GEN_1342;
      end
    end else begin
      buffer_5_info_signed <= _GEN_1342;
    end
    if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          if (3'h5 == checkIndex_2) begin // @[LoadStoreQueue.scala 187:30]
            buffer_5_info_accessWidth <= 2'h0; // @[LoadStoreQueue.scala 187:30]
          end else begin
            buffer_5_info_accessWidth <= _GEN_1350;
          end
        end else begin
          buffer_5_info_accessWidth <= _GEN_1350;
        end
      end else begin
        buffer_5_info_accessWidth <= _GEN_1350;
      end
    end else begin
      buffer_5_info_accessWidth <= _GEN_1350;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_5_addressAndLoadResultTag_threadId <= 1'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_5_addressAndLoadResultTag_threadId <= _GEN_1554;
        end else begin
          buffer_5_addressAndLoadResultTag_threadId <= _GEN_1358;
        end
      end else begin
        buffer_5_addressAndLoadResultTag_threadId <= _GEN_1358;
      end
    end else begin
      buffer_5_addressAndLoadResultTag_threadId <= _GEN_1358;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_5_addressAndLoadResultTag_id <= 4'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_5_addressAndLoadResultTag_id <= _GEN_1562;
        end else begin
          buffer_5_addressAndLoadResultTag_id <= _GEN_1366;
        end
      end else begin
        buffer_5_addressAndLoadResultTag_id <= _GEN_1366;
      end
    end else begin
      buffer_5_addressAndLoadResultTag_id <= _GEN_1366;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_5_address <= 64'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_5_address <= _GEN_1570;
        end else begin
          buffer_5_address <= _GEN_1374;
        end
      end else begin
        buffer_5_address <= _GEN_1374;
      end
    end else begin
      buffer_5_address <= _GEN_1374;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_5_addressValid <= 1'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_5_addressValid <= _GEN_1578;
        end else begin
          buffer_5_addressValid <= _GEN_1382;
        end
      end else begin
        buffer_5_addressValid <= _GEN_1382;
      end
    end else begin
      buffer_5_addressValid <= _GEN_1382;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_5_storeDataTag_threadId <= 1'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_5_storeDataTag_threadId <= _GEN_1586;
        end else begin
          buffer_5_storeDataTag_threadId <= _GEN_1390;
        end
      end else begin
        buffer_5_storeDataTag_threadId <= _GEN_1390;
      end
    end else begin
      buffer_5_storeDataTag_threadId <= _GEN_1390;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_5_storeDataTag_id <= 4'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_5_storeDataTag_id <= _GEN_1594;
        end else begin
          buffer_5_storeDataTag_id <= _GEN_1398;
        end
      end else begin
        buffer_5_storeDataTag_id <= _GEN_1398;
      end
    end else begin
      buffer_5_storeDataTag_id <= _GEN_1398;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_5_storeData <= 64'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_5_storeData <= _GEN_1602;
        end else begin
          buffer_5_storeData <= _GEN_1406;
        end
      end else begin
        buffer_5_storeData <= _GEN_1406;
      end
    end else begin
      buffer_5_storeData <= _GEN_1406;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_5_storeDataValid <= 1'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_5_storeDataValid <= _GEN_1610;
        end else begin
          buffer_5_storeDataValid <= _GEN_1414;
        end
      end else begin
        buffer_5_storeDataValid <= _GEN_1414;
      end
    end else begin
      buffer_5_storeDataValid <= _GEN_1414;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_6_valid <= 1'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_6_valid <= _GEN_1515;
        end else begin
          buffer_6_valid <= _GEN_1319;
        end
      end else begin
        buffer_6_valid <= _GEN_1319;
      end
    end else begin
      buffer_6_valid <= _GEN_1319;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_6_readyReorderSign <= 1'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_6_readyReorderSign <= _GEN_1523;
        end else begin
          buffer_6_readyReorderSign <= _GEN_1327;
        end
      end else begin
        buffer_6_readyReorderSign <= _GEN_1327;
      end
    end else begin
      buffer_6_readyReorderSign <= _GEN_1327;
    end
    if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          if (3'h6 == checkIndex_2) begin // @[LoadStoreQueue.scala 187:30]
            buffer_6_info_accessType <= 1'h0; // @[LoadStoreQueue.scala 187:30]
          end else begin
            buffer_6_info_accessType <= _GEN_1335;
          end
        end else begin
          buffer_6_info_accessType <= _GEN_1335;
        end
      end else begin
        buffer_6_info_accessType <= _GEN_1335;
      end
    end else begin
      buffer_6_info_accessType <= _GEN_1335;
    end
    if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          if (3'h6 == checkIndex_2) begin // @[LoadStoreQueue.scala 187:30]
            buffer_6_info_signed <= 1'h0; // @[LoadStoreQueue.scala 187:30]
          end else begin
            buffer_6_info_signed <= _GEN_1343;
          end
        end else begin
          buffer_6_info_signed <= _GEN_1343;
        end
      end else begin
        buffer_6_info_signed <= _GEN_1343;
      end
    end else begin
      buffer_6_info_signed <= _GEN_1343;
    end
    if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          if (3'h6 == checkIndex_2) begin // @[LoadStoreQueue.scala 187:30]
            buffer_6_info_accessWidth <= 2'h0; // @[LoadStoreQueue.scala 187:30]
          end else begin
            buffer_6_info_accessWidth <= _GEN_1351;
          end
        end else begin
          buffer_6_info_accessWidth <= _GEN_1351;
        end
      end else begin
        buffer_6_info_accessWidth <= _GEN_1351;
      end
    end else begin
      buffer_6_info_accessWidth <= _GEN_1351;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_6_addressAndLoadResultTag_threadId <= 1'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_6_addressAndLoadResultTag_threadId <= _GEN_1555;
        end else begin
          buffer_6_addressAndLoadResultTag_threadId <= _GEN_1359;
        end
      end else begin
        buffer_6_addressAndLoadResultTag_threadId <= _GEN_1359;
      end
    end else begin
      buffer_6_addressAndLoadResultTag_threadId <= _GEN_1359;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_6_addressAndLoadResultTag_id <= 4'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_6_addressAndLoadResultTag_id <= _GEN_1563;
        end else begin
          buffer_6_addressAndLoadResultTag_id <= _GEN_1367;
        end
      end else begin
        buffer_6_addressAndLoadResultTag_id <= _GEN_1367;
      end
    end else begin
      buffer_6_addressAndLoadResultTag_id <= _GEN_1367;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_6_address <= 64'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_6_address <= _GEN_1571;
        end else begin
          buffer_6_address <= _GEN_1375;
        end
      end else begin
        buffer_6_address <= _GEN_1375;
      end
    end else begin
      buffer_6_address <= _GEN_1375;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_6_addressValid <= 1'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_6_addressValid <= _GEN_1579;
        end else begin
          buffer_6_addressValid <= _GEN_1383;
        end
      end else begin
        buffer_6_addressValid <= _GEN_1383;
      end
    end else begin
      buffer_6_addressValid <= _GEN_1383;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_6_storeDataTag_threadId <= 1'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_6_storeDataTag_threadId <= _GEN_1587;
        end else begin
          buffer_6_storeDataTag_threadId <= _GEN_1391;
        end
      end else begin
        buffer_6_storeDataTag_threadId <= _GEN_1391;
      end
    end else begin
      buffer_6_storeDataTag_threadId <= _GEN_1391;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_6_storeDataTag_id <= 4'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_6_storeDataTag_id <= _GEN_1595;
        end else begin
          buffer_6_storeDataTag_id <= _GEN_1399;
        end
      end else begin
        buffer_6_storeDataTag_id <= _GEN_1399;
      end
    end else begin
      buffer_6_storeDataTag_id <= _GEN_1399;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_6_storeData <= 64'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_6_storeData <= _GEN_1603;
        end else begin
          buffer_6_storeData <= _GEN_1407;
        end
      end else begin
        buffer_6_storeData <= _GEN_1407;
      end
    end else begin
      buffer_6_storeData <= _GEN_1407;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_6_storeDataValid <= 1'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_6_storeDataValid <= _GEN_1611;
        end else begin
          buffer_6_storeDataValid <= _GEN_1415;
        end
      end else begin
        buffer_6_storeDataValid <= _GEN_1415;
      end
    end else begin
      buffer_6_storeDataValid <= _GEN_1415;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_7_valid <= 1'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_7_valid <= _GEN_1516;
        end else begin
          buffer_7_valid <= _GEN_1320;
        end
      end else begin
        buffer_7_valid <= _GEN_1320;
      end
    end else begin
      buffer_7_valid <= _GEN_1320;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_7_readyReorderSign <= 1'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_7_readyReorderSign <= _GEN_1524;
        end else begin
          buffer_7_readyReorderSign <= _GEN_1328;
        end
      end else begin
        buffer_7_readyReorderSign <= _GEN_1328;
      end
    end else begin
      buffer_7_readyReorderSign <= _GEN_1328;
    end
    if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          if (3'h7 == checkIndex_2) begin // @[LoadStoreQueue.scala 187:30]
            buffer_7_info_accessType <= 1'h0; // @[LoadStoreQueue.scala 187:30]
          end else begin
            buffer_7_info_accessType <= _GEN_1336;
          end
        end else begin
          buffer_7_info_accessType <= _GEN_1336;
        end
      end else begin
        buffer_7_info_accessType <= _GEN_1336;
      end
    end else begin
      buffer_7_info_accessType <= _GEN_1336;
    end
    if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          if (3'h7 == checkIndex_2) begin // @[LoadStoreQueue.scala 187:30]
            buffer_7_info_signed <= 1'h0; // @[LoadStoreQueue.scala 187:30]
          end else begin
            buffer_7_info_signed <= _GEN_1344;
          end
        end else begin
          buffer_7_info_signed <= _GEN_1344;
        end
      end else begin
        buffer_7_info_signed <= _GEN_1344;
      end
    end else begin
      buffer_7_info_signed <= _GEN_1344;
    end
    if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          if (3'h7 == checkIndex_2) begin // @[LoadStoreQueue.scala 187:30]
            buffer_7_info_accessWidth <= 2'h0; // @[LoadStoreQueue.scala 187:30]
          end else begin
            buffer_7_info_accessWidth <= _GEN_1352;
          end
        end else begin
          buffer_7_info_accessWidth <= _GEN_1352;
        end
      end else begin
        buffer_7_info_accessWidth <= _GEN_1352;
      end
    end else begin
      buffer_7_info_accessWidth <= _GEN_1352;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_7_addressAndLoadResultTag_threadId <= 1'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_7_addressAndLoadResultTag_threadId <= _GEN_1556;
        end else begin
          buffer_7_addressAndLoadResultTag_threadId <= _GEN_1360;
        end
      end else begin
        buffer_7_addressAndLoadResultTag_threadId <= _GEN_1360;
      end
    end else begin
      buffer_7_addressAndLoadResultTag_threadId <= _GEN_1360;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_7_addressAndLoadResultTag_id <= 4'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_7_addressAndLoadResultTag_id <= _GEN_1564;
        end else begin
          buffer_7_addressAndLoadResultTag_id <= _GEN_1368;
        end
      end else begin
        buffer_7_addressAndLoadResultTag_id <= _GEN_1368;
      end
    end else begin
      buffer_7_addressAndLoadResultTag_id <= _GEN_1368;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_7_address <= 64'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_7_address <= _GEN_1572;
        end else begin
          buffer_7_address <= _GEN_1376;
        end
      end else begin
        buffer_7_address <= _GEN_1376;
      end
    end else begin
      buffer_7_address <= _GEN_1376;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_7_addressValid <= 1'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_7_addressValid <= _GEN_1580;
        end else begin
          buffer_7_addressValid <= _GEN_1384;
        end
      end else begin
        buffer_7_addressValid <= _GEN_1384;
      end
    end else begin
      buffer_7_addressValid <= _GEN_1384;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_7_storeDataTag_threadId <= 1'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_7_storeDataTag_threadId <= _GEN_1588;
        end else begin
          buffer_7_storeDataTag_threadId <= _GEN_1392;
        end
      end else begin
        buffer_7_storeDataTag_threadId <= _GEN_1392;
      end
    end else begin
      buffer_7_storeDataTag_threadId <= _GEN_1392;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_7_storeDataTag_id <= 4'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_7_storeDataTag_id <= _GEN_1596;
        end else begin
          buffer_7_storeDataTag_id <= _GEN_1400;
        end
      end else begin
        buffer_7_storeDataTag_id <= _GEN_1400;
      end
    end else begin
      buffer_7_storeDataTag_id <= _GEN_1400;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_7_storeData <= 64'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_7_storeData <= _GEN_1604;
        end else begin
          buffer_7_storeData <= _GEN_1408;
        end
      end else begin
        buffer_7_storeData <= _GEN_1408;
      end
    end else begin
      buffer_7_storeData <= _GEN_1408;
    end
    if (reset) begin // @[LoadStoreQueue.scala 51:23]
      buffer_7_storeDataValid <= 1'h0; // @[LoadStoreQueue.scala 51:23]
    end else if (EntryValid_2) begin // @[LoadStoreQueue.scala 150:36]
      if (checkOk_2 & ~_T_242) begin // @[LoadStoreQueue.scala 181:31]
        if (io_memory_ready) begin // @[LoadStoreQueue.scala 186:31]
          buffer_7_storeDataValid <= _GEN_1612;
        end else begin
          buffer_7_storeDataValid <= _GEN_1416;
        end
      end else begin
        buffer_7_storeDataValid <= _GEN_1416;
      end
    end else begin
      buffer_7_storeDataValid <= _GEN_1416;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  head = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  nextTail = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  buffer_0_valid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  buffer_0_readyReorderSign = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  buffer_0_info_accessType = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  buffer_0_info_signed = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  buffer_0_info_accessWidth = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  buffer_0_addressAndLoadResultTag_threadId = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  buffer_0_addressAndLoadResultTag_id = _RAND_8[3:0];
  _RAND_9 = {2{`RANDOM}};
  buffer_0_address = _RAND_9[63:0];
  _RAND_10 = {1{`RANDOM}};
  buffer_0_addressValid = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  buffer_0_storeDataTag_threadId = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  buffer_0_storeDataTag_id = _RAND_12[3:0];
  _RAND_13 = {2{`RANDOM}};
  buffer_0_storeData = _RAND_13[63:0];
  _RAND_14 = {1{`RANDOM}};
  buffer_0_storeDataValid = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  buffer_1_valid = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  buffer_1_readyReorderSign = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  buffer_1_info_accessType = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  buffer_1_info_signed = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  buffer_1_info_accessWidth = _RAND_19[1:0];
  _RAND_20 = {1{`RANDOM}};
  buffer_1_addressAndLoadResultTag_threadId = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  buffer_1_addressAndLoadResultTag_id = _RAND_21[3:0];
  _RAND_22 = {2{`RANDOM}};
  buffer_1_address = _RAND_22[63:0];
  _RAND_23 = {1{`RANDOM}};
  buffer_1_addressValid = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  buffer_1_storeDataTag_threadId = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  buffer_1_storeDataTag_id = _RAND_25[3:0];
  _RAND_26 = {2{`RANDOM}};
  buffer_1_storeData = _RAND_26[63:0];
  _RAND_27 = {1{`RANDOM}};
  buffer_1_storeDataValid = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  buffer_2_valid = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  buffer_2_readyReorderSign = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  buffer_2_info_accessType = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  buffer_2_info_signed = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  buffer_2_info_accessWidth = _RAND_32[1:0];
  _RAND_33 = {1{`RANDOM}};
  buffer_2_addressAndLoadResultTag_threadId = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  buffer_2_addressAndLoadResultTag_id = _RAND_34[3:0];
  _RAND_35 = {2{`RANDOM}};
  buffer_2_address = _RAND_35[63:0];
  _RAND_36 = {1{`RANDOM}};
  buffer_2_addressValid = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  buffer_2_storeDataTag_threadId = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  buffer_2_storeDataTag_id = _RAND_38[3:0];
  _RAND_39 = {2{`RANDOM}};
  buffer_2_storeData = _RAND_39[63:0];
  _RAND_40 = {1{`RANDOM}};
  buffer_2_storeDataValid = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  buffer_3_valid = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  buffer_3_readyReorderSign = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  buffer_3_info_accessType = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  buffer_3_info_signed = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  buffer_3_info_accessWidth = _RAND_45[1:0];
  _RAND_46 = {1{`RANDOM}};
  buffer_3_addressAndLoadResultTag_threadId = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  buffer_3_addressAndLoadResultTag_id = _RAND_47[3:0];
  _RAND_48 = {2{`RANDOM}};
  buffer_3_address = _RAND_48[63:0];
  _RAND_49 = {1{`RANDOM}};
  buffer_3_addressValid = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  buffer_3_storeDataTag_threadId = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  buffer_3_storeDataTag_id = _RAND_51[3:0];
  _RAND_52 = {2{`RANDOM}};
  buffer_3_storeData = _RAND_52[63:0];
  _RAND_53 = {1{`RANDOM}};
  buffer_3_storeDataValid = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  buffer_4_valid = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  buffer_4_readyReorderSign = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  buffer_4_info_accessType = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  buffer_4_info_signed = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  buffer_4_info_accessWidth = _RAND_58[1:0];
  _RAND_59 = {1{`RANDOM}};
  buffer_4_addressAndLoadResultTag_threadId = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  buffer_4_addressAndLoadResultTag_id = _RAND_60[3:0];
  _RAND_61 = {2{`RANDOM}};
  buffer_4_address = _RAND_61[63:0];
  _RAND_62 = {1{`RANDOM}};
  buffer_4_addressValid = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  buffer_4_storeDataTag_threadId = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  buffer_4_storeDataTag_id = _RAND_64[3:0];
  _RAND_65 = {2{`RANDOM}};
  buffer_4_storeData = _RAND_65[63:0];
  _RAND_66 = {1{`RANDOM}};
  buffer_4_storeDataValid = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  buffer_5_valid = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  buffer_5_readyReorderSign = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  buffer_5_info_accessType = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  buffer_5_info_signed = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  buffer_5_info_accessWidth = _RAND_71[1:0];
  _RAND_72 = {1{`RANDOM}};
  buffer_5_addressAndLoadResultTag_threadId = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  buffer_5_addressAndLoadResultTag_id = _RAND_73[3:0];
  _RAND_74 = {2{`RANDOM}};
  buffer_5_address = _RAND_74[63:0];
  _RAND_75 = {1{`RANDOM}};
  buffer_5_addressValid = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  buffer_5_storeDataTag_threadId = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  buffer_5_storeDataTag_id = _RAND_77[3:0];
  _RAND_78 = {2{`RANDOM}};
  buffer_5_storeData = _RAND_78[63:0];
  _RAND_79 = {1{`RANDOM}};
  buffer_5_storeDataValid = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  buffer_6_valid = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  buffer_6_readyReorderSign = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  buffer_6_info_accessType = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  buffer_6_info_signed = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  buffer_6_info_accessWidth = _RAND_84[1:0];
  _RAND_85 = {1{`RANDOM}};
  buffer_6_addressAndLoadResultTag_threadId = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  buffer_6_addressAndLoadResultTag_id = _RAND_86[3:0];
  _RAND_87 = {2{`RANDOM}};
  buffer_6_address = _RAND_87[63:0];
  _RAND_88 = {1{`RANDOM}};
  buffer_6_addressValid = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  buffer_6_storeDataTag_threadId = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  buffer_6_storeDataTag_id = _RAND_90[3:0];
  _RAND_91 = {2{`RANDOM}};
  buffer_6_storeData = _RAND_91[63:0];
  _RAND_92 = {1{`RANDOM}};
  buffer_6_storeDataValid = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  buffer_7_valid = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  buffer_7_readyReorderSign = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  buffer_7_info_accessType = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  buffer_7_info_signed = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  buffer_7_info_accessWidth = _RAND_97[1:0];
  _RAND_98 = {1{`RANDOM}};
  buffer_7_addressAndLoadResultTag_threadId = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  buffer_7_addressAndLoadResultTag_id = _RAND_99[3:0];
  _RAND_100 = {2{`RANDOM}};
  buffer_7_address = _RAND_100[63:0];
  _RAND_101 = {1{`RANDOM}};
  buffer_7_addressValid = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  buffer_7_storeDataTag_threadId = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  buffer_7_storeDataTag_id = _RAND_103[3:0];
  _RAND_104 = {2{`RANDOM}};
  buffer_7_storeData = _RAND_104[63:0];
  _RAND_105 = {1{`RANDOM}};
  buffer_7_storeDataValid = _RAND_105[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module B4RRArbiter(
  input         clock,
  input         reset,
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [63:0] io_in_0_bits_address,
  input         io_in_0_bits_tag_threadId,
  input  [3:0]  io_in_0_bits_tag_id,
  input  [63:0] io_in_0_bits_data,
  input         io_in_0_bits_accessInfo_accessType,
  input         io_in_0_bits_accessInfo_signed,
  input  [1:0]  io_in_0_bits_accessInfo_accessWidth,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [63:0] io_in_1_bits_address,
  input         io_in_1_bits_tag_threadId,
  input  [3:0]  io_in_1_bits_tag_id,
  input  [63:0] io_in_1_bits_data,
  input         io_in_1_bits_accessInfo_accessType,
  input         io_in_1_bits_accessInfo_signed,
  input  [1:0]  io_in_1_bits_accessInfo_accessWidth,
  input         io_out_ready,
  output        io_out_valid,
  output [63:0] io_out_bits_address,
  output        io_out_bits_tag_threadId,
  output [3:0]  io_out_bits_tag_id,
  output [63:0] io_out_bits_data,
  output        io_out_bits_accessInfo_accessType,
  output        io_out_bits_accessInfo_signed,
  output [1:0]  io_out_bits_accessInfo_accessWidth,
  output        io_chosen
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  _ctrl_validMask_grantMask_lastGrant_T = io_out_ready & io_out_valid; // @[Decoupled.scala 51:35]
  reg  lastGrant; // @[Reg.scala 35:20]
  wire  grantMask_1 = 1'h1 > lastGrant; // @[Arbitar.scala 89:49]
  wire  validMask_1 = io_in_1_valid & grantMask_1; // @[Arbitar.scala 91:57]
  wire  ctrl_2 = ~validMask_1; // @[Arbitar.scala 44:78]
  wire  ctrl_3 = ~(validMask_1 | io_in_0_valid); // @[Arbitar.scala 44:78]
  wire  _T_3 = grantMask_1 | ctrl_3; // @[Arbitar.scala 97:50]
  wire  _GEN_17 = io_in_0_valid ? 1'h0 : 1'h1; // @[Arbitar.scala 102:{26,35} 100:41]
  assign io_in_0_ready = ctrl_2 & io_out_ready; // @[Arbitar.scala 78:21]
  assign io_in_1_ready = _T_3 & io_out_ready; // @[Arbitar.scala 78:21]
  assign io_out_valid = io_chosen ? io_in_1_valid : io_in_0_valid; // @[Arbitar.scala 59:{16,16}]
  assign io_out_bits_address = io_chosen ? io_in_1_bits_address : io_in_0_bits_address; // @[Arbitar.scala 60:{15,15}]
  assign io_out_bits_tag_threadId = io_chosen ? io_in_1_bits_tag_threadId : io_in_0_bits_tag_threadId; // @[Arbitar.scala 60:{15,15}]
  assign io_out_bits_tag_id = io_chosen ? io_in_1_bits_tag_id : io_in_0_bits_tag_id; // @[Arbitar.scala 60:{15,15}]
  assign io_out_bits_data = io_chosen ? io_in_1_bits_data : io_in_0_bits_data; // @[Arbitar.scala 60:{15,15}]
  assign io_out_bits_accessInfo_accessType = io_chosen ? io_in_1_bits_accessInfo_accessType :
    io_in_0_bits_accessInfo_accessType; // @[Arbitar.scala 60:{15,15}]
  assign io_out_bits_accessInfo_signed = io_chosen ? io_in_1_bits_accessInfo_signed : io_in_0_bits_accessInfo_signed; // @[Arbitar.scala 60:{15,15}]
  assign io_out_bits_accessInfo_accessWidth = io_chosen ? io_in_1_bits_accessInfo_accessWidth :
    io_in_0_bits_accessInfo_accessWidth; // @[Arbitar.scala 60:{15,15}]
  assign io_chosen = validMask_1 | _GEN_17; // @[Arbitar.scala 104:{24,33}]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 35:20]
      lastGrant <= 1'h0; // @[Reg.scala 35:20]
    end else if (_ctrl_validMask_grantMask_lastGrant_T) begin // @[Reg.scala 36:18]
      lastGrant <= io_chosen; // @[Reg.scala 36:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  lastGrant = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [63:0] io_enq_bits_address,
  input         io_enq_bits_tag_threadId,
  input  [3:0]  io_enq_bits_tag_id,
  input  [63:0] io_enq_bits_data,
  input         io_enq_bits_accessInfo_accessType,
  input         io_enq_bits_accessInfo_signed,
  input  [1:0]  io_enq_bits_accessInfo_accessWidth,
  input         io_deq_ready,
  output        io_deq_valid,
  output [63:0] io_deq_bits_address,
  output        io_deq_bits_tag_threadId,
  output [3:0]  io_deq_bits_tag_id,
  output [63:0] io_deq_bits_data,
  output        io_deq_bits_accessInfo_accessType,
  output        io_deq_bits_accessInfo_signed,
  output [1:0]  io_deq_bits_accessInfo_accessWidth
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_6;
  reg [63:0] _RAND_9;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_18;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] ram_address [0:7]; // @[Decoupled.scala 273:44]
  wire  ram_address_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:44]
  wire [2:0] ram_address_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:44]
  wire [63:0] ram_address_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:44]
  wire [63:0] ram_address_MPORT_data; // @[Decoupled.scala 273:44]
  wire [2:0] ram_address_MPORT_addr; // @[Decoupled.scala 273:44]
  wire  ram_address_MPORT_mask; // @[Decoupled.scala 273:44]
  wire  ram_address_MPORT_en; // @[Decoupled.scala 273:44]
  reg  ram_address_io_deq_bits_MPORT_en_pipe_0;
  reg [2:0] ram_address_io_deq_bits_MPORT_addr_pipe_0;
  reg  ram_tag_threadId [0:7]; // @[Decoupled.scala 273:44]
  wire  ram_tag_threadId_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:44]
  wire [2:0] ram_tag_threadId_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:44]
  wire  ram_tag_threadId_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:44]
  wire  ram_tag_threadId_MPORT_data; // @[Decoupled.scala 273:44]
  wire [2:0] ram_tag_threadId_MPORT_addr; // @[Decoupled.scala 273:44]
  wire  ram_tag_threadId_MPORT_mask; // @[Decoupled.scala 273:44]
  wire  ram_tag_threadId_MPORT_en; // @[Decoupled.scala 273:44]
  reg  ram_tag_threadId_io_deq_bits_MPORT_en_pipe_0;
  reg [2:0] ram_tag_threadId_io_deq_bits_MPORT_addr_pipe_0;
  reg [3:0] ram_tag_id [0:7]; // @[Decoupled.scala 273:44]
  wire  ram_tag_id_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:44]
  wire [2:0] ram_tag_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:44]
  wire [3:0] ram_tag_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:44]
  wire [3:0] ram_tag_id_MPORT_data; // @[Decoupled.scala 273:44]
  wire [2:0] ram_tag_id_MPORT_addr; // @[Decoupled.scala 273:44]
  wire  ram_tag_id_MPORT_mask; // @[Decoupled.scala 273:44]
  wire  ram_tag_id_MPORT_en; // @[Decoupled.scala 273:44]
  reg  ram_tag_id_io_deq_bits_MPORT_en_pipe_0;
  reg [2:0] ram_tag_id_io_deq_bits_MPORT_addr_pipe_0;
  reg [63:0] ram_data [0:7]; // @[Decoupled.scala 273:44]
  wire  ram_data_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:44]
  wire [2:0] ram_data_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:44]
  wire [63:0] ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:44]
  wire [63:0] ram_data_MPORT_data; // @[Decoupled.scala 273:44]
  wire [2:0] ram_data_MPORT_addr; // @[Decoupled.scala 273:44]
  wire  ram_data_MPORT_mask; // @[Decoupled.scala 273:44]
  wire  ram_data_MPORT_en; // @[Decoupled.scala 273:44]
  reg  ram_data_io_deq_bits_MPORT_en_pipe_0;
  reg [2:0] ram_data_io_deq_bits_MPORT_addr_pipe_0;
  reg  ram_accessInfo_accessType [0:7]; // @[Decoupled.scala 273:44]
  wire  ram_accessInfo_accessType_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:44]
  wire [2:0] ram_accessInfo_accessType_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:44]
  wire  ram_accessInfo_accessType_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:44]
  wire  ram_accessInfo_accessType_MPORT_data; // @[Decoupled.scala 273:44]
  wire [2:0] ram_accessInfo_accessType_MPORT_addr; // @[Decoupled.scala 273:44]
  wire  ram_accessInfo_accessType_MPORT_mask; // @[Decoupled.scala 273:44]
  wire  ram_accessInfo_accessType_MPORT_en; // @[Decoupled.scala 273:44]
  reg  ram_accessInfo_accessType_io_deq_bits_MPORT_en_pipe_0;
  reg [2:0] ram_accessInfo_accessType_io_deq_bits_MPORT_addr_pipe_0;
  reg  ram_accessInfo_signed [0:7]; // @[Decoupled.scala 273:44]
  wire  ram_accessInfo_signed_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:44]
  wire [2:0] ram_accessInfo_signed_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:44]
  wire  ram_accessInfo_signed_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:44]
  wire  ram_accessInfo_signed_MPORT_data; // @[Decoupled.scala 273:44]
  wire [2:0] ram_accessInfo_signed_MPORT_addr; // @[Decoupled.scala 273:44]
  wire  ram_accessInfo_signed_MPORT_mask; // @[Decoupled.scala 273:44]
  wire  ram_accessInfo_signed_MPORT_en; // @[Decoupled.scala 273:44]
  reg  ram_accessInfo_signed_io_deq_bits_MPORT_en_pipe_0;
  reg [2:0] ram_accessInfo_signed_io_deq_bits_MPORT_addr_pipe_0;
  reg [1:0] ram_accessInfo_accessWidth [0:7]; // @[Decoupled.scala 273:44]
  wire  ram_accessInfo_accessWidth_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:44]
  wire [2:0] ram_accessInfo_accessWidth_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:44]
  wire [1:0] ram_accessInfo_accessWidth_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:44]
  wire [1:0] ram_accessInfo_accessWidth_MPORT_data; // @[Decoupled.scala 273:44]
  wire [2:0] ram_accessInfo_accessWidth_MPORT_addr; // @[Decoupled.scala 273:44]
  wire  ram_accessInfo_accessWidth_MPORT_mask; // @[Decoupled.scala 273:44]
  wire  ram_accessInfo_accessWidth_MPORT_en; // @[Decoupled.scala 273:44]
  reg  ram_accessInfo_accessWidth_io_deq_bits_MPORT_en_pipe_0;
  reg [2:0] ram_accessInfo_accessWidth_io_deq_bits_MPORT_addr_pipe_0;
  reg [2:0] enq_ptr_value; // @[Counter.scala 61:40]
  reg [2:0] deq_ptr_value; // @[Counter.scala 61:40]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 277:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 278:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 279:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _value_T_1 = enq_ptr_value + 3'h1; // @[Counter.scala 77:24]
  wire [2:0] _value_T_3 = deq_ptr_value + 3'h1; // @[Counter.scala 77:24]
  wire [3:0] _deq_ptr_next_T_1 = 4'h8 - 4'h1; // @[Decoupled.scala 306:57]
  wire [3:0] _GEN_21 = {{1'd0}, deq_ptr_value}; // @[Decoupled.scala 306:42]
  assign ram_address_io_deq_bits_MPORT_en = ram_address_io_deq_bits_MPORT_en_pipe_0;
  assign ram_address_io_deq_bits_MPORT_addr = ram_address_io_deq_bits_MPORT_addr_pipe_0;
  assign ram_address_io_deq_bits_MPORT_data = ram_address[ram_address_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:44]
  assign ram_address_MPORT_data = io_enq_bits_address;
  assign ram_address_MPORT_addr = enq_ptr_value;
  assign ram_address_MPORT_mask = 1'h1;
  assign ram_address_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_tag_threadId_io_deq_bits_MPORT_en = ram_tag_threadId_io_deq_bits_MPORT_en_pipe_0;
  assign ram_tag_threadId_io_deq_bits_MPORT_addr = ram_tag_threadId_io_deq_bits_MPORT_addr_pipe_0;
  assign ram_tag_threadId_io_deq_bits_MPORT_data = ram_tag_threadId[ram_tag_threadId_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:44]
  assign ram_tag_threadId_MPORT_data = io_enq_bits_tag_threadId;
  assign ram_tag_threadId_MPORT_addr = enq_ptr_value;
  assign ram_tag_threadId_MPORT_mask = 1'h1;
  assign ram_tag_threadId_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_tag_id_io_deq_bits_MPORT_en = ram_tag_id_io_deq_bits_MPORT_en_pipe_0;
  assign ram_tag_id_io_deq_bits_MPORT_addr = ram_tag_id_io_deq_bits_MPORT_addr_pipe_0;
  assign ram_tag_id_io_deq_bits_MPORT_data = ram_tag_id[ram_tag_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:44]
  assign ram_tag_id_MPORT_data = io_enq_bits_tag_id;
  assign ram_tag_id_MPORT_addr = enq_ptr_value;
  assign ram_tag_id_MPORT_mask = 1'h1;
  assign ram_tag_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_data_io_deq_bits_MPORT_en = ram_data_io_deq_bits_MPORT_en_pipe_0;
  assign ram_data_io_deq_bits_MPORT_addr = ram_data_io_deq_bits_MPORT_addr_pipe_0;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:44]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = enq_ptr_value;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_accessInfo_accessType_io_deq_bits_MPORT_en = ram_accessInfo_accessType_io_deq_bits_MPORT_en_pipe_0;
  assign ram_accessInfo_accessType_io_deq_bits_MPORT_addr = ram_accessInfo_accessType_io_deq_bits_MPORT_addr_pipe_0;
  assign ram_accessInfo_accessType_io_deq_bits_MPORT_data =
    ram_accessInfo_accessType[ram_accessInfo_accessType_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:44]
  assign ram_accessInfo_accessType_MPORT_data = io_enq_bits_accessInfo_accessType;
  assign ram_accessInfo_accessType_MPORT_addr = enq_ptr_value;
  assign ram_accessInfo_accessType_MPORT_mask = 1'h1;
  assign ram_accessInfo_accessType_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_accessInfo_signed_io_deq_bits_MPORT_en = ram_accessInfo_signed_io_deq_bits_MPORT_en_pipe_0;
  assign ram_accessInfo_signed_io_deq_bits_MPORT_addr = ram_accessInfo_signed_io_deq_bits_MPORT_addr_pipe_0;
  assign ram_accessInfo_signed_io_deq_bits_MPORT_data =
    ram_accessInfo_signed[ram_accessInfo_signed_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:44]
  assign ram_accessInfo_signed_MPORT_data = io_enq_bits_accessInfo_signed;
  assign ram_accessInfo_signed_MPORT_addr = enq_ptr_value;
  assign ram_accessInfo_signed_MPORT_mask = 1'h1;
  assign ram_accessInfo_signed_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_accessInfo_accessWidth_io_deq_bits_MPORT_en = ram_accessInfo_accessWidth_io_deq_bits_MPORT_en_pipe_0;
  assign ram_accessInfo_accessWidth_io_deq_bits_MPORT_addr = ram_accessInfo_accessWidth_io_deq_bits_MPORT_addr_pipe_0;
  assign ram_accessInfo_accessWidth_io_deq_bits_MPORT_data =
    ram_accessInfo_accessWidth[ram_accessInfo_accessWidth_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:44]
  assign ram_accessInfo_accessWidth_MPORT_data = io_enq_bits_accessInfo_accessWidth;
  assign ram_accessInfo_accessWidth_MPORT_addr = enq_ptr_value;
  assign ram_accessInfo_accessWidth_MPORT_mask = 1'h1;
  assign ram_accessInfo_accessWidth_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 303:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 302:19]
  assign io_deq_bits_address = ram_address_io_deq_bits_MPORT_data; // @[Decoupled.scala 308:17]
  assign io_deq_bits_tag_threadId = ram_tag_threadId_io_deq_bits_MPORT_data; // @[Decoupled.scala 308:17]
  assign io_deq_bits_tag_id = ram_tag_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 308:17]
  assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 308:17]
  assign io_deq_bits_accessInfo_accessType = ram_accessInfo_accessType_io_deq_bits_MPORT_data; // @[Decoupled.scala 308:17]
  assign io_deq_bits_accessInfo_signed = ram_accessInfo_signed_io_deq_bits_MPORT_data; // @[Decoupled.scala 308:17]
  assign io_deq_bits_accessInfo_accessWidth = ram_accessInfo_accessWidth_io_deq_bits_MPORT_data; // @[Decoupled.scala 308:17]
  always @(posedge clock) begin
    if (ram_address_MPORT_en & ram_address_MPORT_mask) begin
      ram_address[ram_address_MPORT_addr] <= ram_address_MPORT_data; // @[Decoupled.scala 273:44]
    end
    ram_address_io_deq_bits_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (do_deq) begin
        if (_GEN_21 == _deq_ptr_next_T_1) begin // @[Decoupled.scala 306:27]
          ram_address_io_deq_bits_MPORT_addr_pipe_0 <= 3'h0;
        end else begin
          ram_address_io_deq_bits_MPORT_addr_pipe_0 <= _value_T_3;
        end
      end else begin
        ram_address_io_deq_bits_MPORT_addr_pipe_0 <= deq_ptr_value;
      end
    end
    if (ram_tag_threadId_MPORT_en & ram_tag_threadId_MPORT_mask) begin
      ram_tag_threadId[ram_tag_threadId_MPORT_addr] <= ram_tag_threadId_MPORT_data; // @[Decoupled.scala 273:44]
    end
    ram_tag_threadId_io_deq_bits_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (do_deq) begin
        if (_GEN_21 == _deq_ptr_next_T_1) begin // @[Decoupled.scala 306:27]
          ram_tag_threadId_io_deq_bits_MPORT_addr_pipe_0 <= 3'h0;
        end else begin
          ram_tag_threadId_io_deq_bits_MPORT_addr_pipe_0 <= _value_T_3;
        end
      end else begin
        ram_tag_threadId_io_deq_bits_MPORT_addr_pipe_0 <= deq_ptr_value;
      end
    end
    if (ram_tag_id_MPORT_en & ram_tag_id_MPORT_mask) begin
      ram_tag_id[ram_tag_id_MPORT_addr] <= ram_tag_id_MPORT_data; // @[Decoupled.scala 273:44]
    end
    ram_tag_id_io_deq_bits_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (do_deq) begin
        if (_GEN_21 == _deq_ptr_next_T_1) begin // @[Decoupled.scala 306:27]
          ram_tag_id_io_deq_bits_MPORT_addr_pipe_0 <= 3'h0;
        end else begin
          ram_tag_id_io_deq_bits_MPORT_addr_pipe_0 <= _value_T_3;
        end
      end else begin
        ram_tag_id_io_deq_bits_MPORT_addr_pipe_0 <= deq_ptr_value;
      end
    end
    if (ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[Decoupled.scala 273:44]
    end
    ram_data_io_deq_bits_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (do_deq) begin
        if (_GEN_21 == _deq_ptr_next_T_1) begin // @[Decoupled.scala 306:27]
          ram_data_io_deq_bits_MPORT_addr_pipe_0 <= 3'h0;
        end else begin
          ram_data_io_deq_bits_MPORT_addr_pipe_0 <= _value_T_3;
        end
      end else begin
        ram_data_io_deq_bits_MPORT_addr_pipe_0 <= deq_ptr_value;
      end
    end
    if (ram_accessInfo_accessType_MPORT_en & ram_accessInfo_accessType_MPORT_mask) begin
      ram_accessInfo_accessType[ram_accessInfo_accessType_MPORT_addr] <= ram_accessInfo_accessType_MPORT_data; // @[Decoupled.scala 273:44]
    end
    ram_accessInfo_accessType_io_deq_bits_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (do_deq) begin
        if (_GEN_21 == _deq_ptr_next_T_1) begin // @[Decoupled.scala 306:27]
          ram_accessInfo_accessType_io_deq_bits_MPORT_addr_pipe_0 <= 3'h0;
        end else begin
          ram_accessInfo_accessType_io_deq_bits_MPORT_addr_pipe_0 <= _value_T_3;
        end
      end else begin
        ram_accessInfo_accessType_io_deq_bits_MPORT_addr_pipe_0 <= deq_ptr_value;
      end
    end
    if (ram_accessInfo_signed_MPORT_en & ram_accessInfo_signed_MPORT_mask) begin
      ram_accessInfo_signed[ram_accessInfo_signed_MPORT_addr] <= ram_accessInfo_signed_MPORT_data; // @[Decoupled.scala 273:44]
    end
    ram_accessInfo_signed_io_deq_bits_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (do_deq) begin
        if (_GEN_21 == _deq_ptr_next_T_1) begin // @[Decoupled.scala 306:27]
          ram_accessInfo_signed_io_deq_bits_MPORT_addr_pipe_0 <= 3'h0;
        end else begin
          ram_accessInfo_signed_io_deq_bits_MPORT_addr_pipe_0 <= _value_T_3;
        end
      end else begin
        ram_accessInfo_signed_io_deq_bits_MPORT_addr_pipe_0 <= deq_ptr_value;
      end
    end
    if (ram_accessInfo_accessWidth_MPORT_en & ram_accessInfo_accessWidth_MPORT_mask) begin
      ram_accessInfo_accessWidth[ram_accessInfo_accessWidth_MPORT_addr] <= ram_accessInfo_accessWidth_MPORT_data; // @[Decoupled.scala 273:44]
    end
    ram_accessInfo_accessWidth_io_deq_bits_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (do_deq) begin
        if (_GEN_21 == _deq_ptr_next_T_1) begin // @[Decoupled.scala 306:27]
          ram_accessInfo_accessWidth_io_deq_bits_MPORT_addr_pipe_0 <= 3'h0;
        end else begin
          ram_accessInfo_accessWidth_io_deq_bits_MPORT_addr_pipe_0 <= _value_T_3;
        end
      end else begin
        ram_accessInfo_accessWidth_io_deq_bits_MPORT_addr_pipe_0 <= deq_ptr_value;
      end
    end
    if (reset) begin // @[Counter.scala 61:40]
      enq_ptr_value <= 3'h0; // @[Counter.scala 61:40]
    end else if (do_enq) begin // @[Decoupled.scala 286:16]
      enq_ptr_value <= _value_T_1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      deq_ptr_value <= 3'h0; // @[Counter.scala 61:40]
    end else if (do_deq) begin // @[Decoupled.scala 290:16]
      deq_ptr_value <= _value_T_3; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      maybe_full <= do_enq; // @[Decoupled.scala 294:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_address[initvar] = _RAND_0[63:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_tag_threadId[initvar] = _RAND_3[0:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_tag_id[initvar] = _RAND_6[3:0];
  _RAND_9 = {2{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_data[initvar] = _RAND_9[63:0];
  _RAND_12 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_accessInfo_accessType[initvar] = _RAND_12[0:0];
  _RAND_15 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_accessInfo_signed[initvar] = _RAND_15[0:0];
  _RAND_18 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_accessInfo_accessWidth[initvar] = _RAND_18[1:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_address_io_deq_bits_MPORT_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  ram_address_io_deq_bits_MPORT_addr_pipe_0 = _RAND_2[2:0];
  _RAND_4 = {1{`RANDOM}};
  ram_tag_threadId_io_deq_bits_MPORT_en_pipe_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  ram_tag_threadId_io_deq_bits_MPORT_addr_pipe_0 = _RAND_5[2:0];
  _RAND_7 = {1{`RANDOM}};
  ram_tag_id_io_deq_bits_MPORT_en_pipe_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  ram_tag_id_io_deq_bits_MPORT_addr_pipe_0 = _RAND_8[2:0];
  _RAND_10 = {1{`RANDOM}};
  ram_data_io_deq_bits_MPORT_en_pipe_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  ram_data_io_deq_bits_MPORT_addr_pipe_0 = _RAND_11[2:0];
  _RAND_13 = {1{`RANDOM}};
  ram_accessInfo_accessType_io_deq_bits_MPORT_en_pipe_0 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  ram_accessInfo_accessType_io_deq_bits_MPORT_addr_pipe_0 = _RAND_14[2:0];
  _RAND_16 = {1{`RANDOM}};
  ram_accessInfo_signed_io_deq_bits_MPORT_en_pipe_0 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  ram_accessInfo_signed_io_deq_bits_MPORT_addr_pipe_0 = _RAND_17[2:0];
  _RAND_19 = {1{`RANDOM}};
  ram_accessInfo_accessWidth_io_deq_bits_MPORT_en_pipe_0 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  ram_accessInfo_accessWidth_io_deq_bits_MPORT_addr_pipe_0 = _RAND_20[2:0];
  _RAND_21 = {1{`RANDOM}};
  enq_ptr_value = _RAND_21[2:0];
  _RAND_22 = {1{`RANDOM}};
  deq_ptr_value = _RAND_22[2:0];
  _RAND_23 = {1{`RANDOM}};
  maybe_full = _RAND_23[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module FIFO(
  input         clock,
  input         reset,
  output        input_ready,
  input         input_valid,
  input  [63:0] input_bits_address,
  input         input_bits_tag_threadId,
  input  [3:0]  input_bits_tag_id,
  input  [63:0] input_bits_data,
  input         input_bits_accessInfo_accessType,
  input         input_bits_accessInfo_signed,
  input  [1:0]  input_bits_accessInfo_accessWidth,
  input         output_ready,
  output [63:0] output_bits_address,
  output        output_bits_tag_threadId,
  output [3:0]  output_bits_tag_id,
  output [63:0] output_bits_data,
  output        output_bits_accessInfo_accessType,
  output        output_bits_accessInfo_signed,
  output [1:0]  output_bits_accessInfo_accessWidth,
  output        empty
);
  wire  queue_clock; // @[FIFO.scala 16:29]
  wire  queue_reset; // @[FIFO.scala 16:29]
  wire  queue_io_enq_ready; // @[FIFO.scala 16:29]
  wire  queue_io_enq_valid; // @[FIFO.scala 16:29]
  wire [63:0] queue_io_enq_bits_address; // @[FIFO.scala 16:29]
  wire  queue_io_enq_bits_tag_threadId; // @[FIFO.scala 16:29]
  wire [3:0] queue_io_enq_bits_tag_id; // @[FIFO.scala 16:29]
  wire [63:0] queue_io_enq_bits_data; // @[FIFO.scala 16:29]
  wire  queue_io_enq_bits_accessInfo_accessType; // @[FIFO.scala 16:29]
  wire  queue_io_enq_bits_accessInfo_signed; // @[FIFO.scala 16:29]
  wire [1:0] queue_io_enq_bits_accessInfo_accessWidth; // @[FIFO.scala 16:29]
  wire  queue_io_deq_ready; // @[FIFO.scala 16:29]
  wire  queue_io_deq_valid; // @[FIFO.scala 16:29]
  wire [63:0] queue_io_deq_bits_address; // @[FIFO.scala 16:29]
  wire  queue_io_deq_bits_tag_threadId; // @[FIFO.scala 16:29]
  wire [3:0] queue_io_deq_bits_tag_id; // @[FIFO.scala 16:29]
  wire [63:0] queue_io_deq_bits_data; // @[FIFO.scala 16:29]
  wire  queue_io_deq_bits_accessInfo_accessType; // @[FIFO.scala 16:29]
  wire  queue_io_deq_bits_accessInfo_signed; // @[FIFO.scala 16:29]
  wire [1:0] queue_io_deq_bits_accessInfo_accessWidth; // @[FIFO.scala 16:29]
  Queue queue ( // @[FIFO.scala 16:29]
    .clock(queue_clock),
    .reset(queue_reset),
    .io_enq_ready(queue_io_enq_ready),
    .io_enq_valid(queue_io_enq_valid),
    .io_enq_bits_address(queue_io_enq_bits_address),
    .io_enq_bits_tag_threadId(queue_io_enq_bits_tag_threadId),
    .io_enq_bits_tag_id(queue_io_enq_bits_tag_id),
    .io_enq_bits_data(queue_io_enq_bits_data),
    .io_enq_bits_accessInfo_accessType(queue_io_enq_bits_accessInfo_accessType),
    .io_enq_bits_accessInfo_signed(queue_io_enq_bits_accessInfo_signed),
    .io_enq_bits_accessInfo_accessWidth(queue_io_enq_bits_accessInfo_accessWidth),
    .io_deq_ready(queue_io_deq_ready),
    .io_deq_valid(queue_io_deq_valid),
    .io_deq_bits_address(queue_io_deq_bits_address),
    .io_deq_bits_tag_threadId(queue_io_deq_bits_tag_threadId),
    .io_deq_bits_tag_id(queue_io_deq_bits_tag_id),
    .io_deq_bits_data(queue_io_deq_bits_data),
    .io_deq_bits_accessInfo_accessType(queue_io_deq_bits_accessInfo_accessType),
    .io_deq_bits_accessInfo_signed(queue_io_deq_bits_accessInfo_signed),
    .io_deq_bits_accessInfo_accessWidth(queue_io_deq_bits_accessInfo_accessWidth)
  );
  assign input_ready = queue_io_enq_ready; // @[FIFO.scala 19:16]
  assign output_bits_address = queue_io_deq_bits_address; // @[FIFO.scala 20:10]
  assign output_bits_tag_threadId = queue_io_deq_bits_tag_threadId; // @[FIFO.scala 20:10]
  assign output_bits_tag_id = queue_io_deq_bits_tag_id; // @[FIFO.scala 20:10]
  assign output_bits_data = queue_io_deq_bits_data; // @[FIFO.scala 20:10]
  assign output_bits_accessInfo_accessType = queue_io_deq_bits_accessInfo_accessType; // @[FIFO.scala 20:10]
  assign output_bits_accessInfo_signed = queue_io_deq_bits_accessInfo_signed; // @[FIFO.scala 20:10]
  assign output_bits_accessInfo_accessWidth = queue_io_deq_bits_accessInfo_accessWidth; // @[FIFO.scala 20:10]
  assign empty = ~queue_io_deq_valid; // @[FIFO.scala 22:12]
  assign queue_clock = clock;
  assign queue_reset = reset;
  assign queue_io_enq_valid = input_valid; // @[FIFO.scala 19:16]
  assign queue_io_enq_bits_address = input_bits_address; // @[FIFO.scala 19:16]
  assign queue_io_enq_bits_tag_threadId = input_bits_tag_threadId; // @[FIFO.scala 19:16]
  assign queue_io_enq_bits_tag_id = input_bits_tag_id; // @[FIFO.scala 19:16]
  assign queue_io_enq_bits_data = input_bits_data; // @[FIFO.scala 19:16]
  assign queue_io_enq_bits_accessInfo_accessType = input_bits_accessInfo_accessType; // @[FIFO.scala 19:16]
  assign queue_io_enq_bits_accessInfo_signed = input_bits_accessInfo_signed; // @[FIFO.scala 19:16]
  assign queue_io_enq_bits_accessInfo_accessWidth = input_bits_accessInfo_accessWidth; // @[FIFO.scala 19:16]
  assign queue_io_deq_ready = output_ready; // @[FIFO.scala 20:10]
endmodule
module DataMemoryBuffer(
  input         clock,
  input         reset,
  output        io_dataIn_0_ready,
  input         io_dataIn_0_valid,
  input  [63:0] io_dataIn_0_bits_address,
  input         io_dataIn_0_bits_tag_threadId,
  input  [3:0]  io_dataIn_0_bits_tag_id,
  input  [63:0] io_dataIn_0_bits_data,
  input         io_dataIn_0_bits_accessInfo_accessType,
  input         io_dataIn_0_bits_accessInfo_signed,
  input  [1:0]  io_dataIn_0_bits_accessInfo_accessWidth,
  output        io_dataIn_1_ready,
  input         io_dataIn_1_valid,
  input  [63:0] io_dataIn_1_bits_address,
  input         io_dataIn_1_bits_tag_threadId,
  input  [3:0]  io_dataIn_1_bits_tag_id,
  input  [63:0] io_dataIn_1_bits_data,
  input         io_dataIn_1_bits_accessInfo_accessType,
  input         io_dataIn_1_bits_accessInfo_signed,
  input  [1:0]  io_dataIn_1_bits_accessInfo_accessWidth,
  input         io_dataReadRequest_ready,
  output        io_dataReadRequest_valid,
  output [63:0] io_dataReadRequest_bits_address,
  output [1:0]  io_dataReadRequest_bits_size,
  output        io_dataReadRequest_bits_signed,
  output        io_dataReadRequest_bits_outputTag_threadId,
  output [3:0]  io_dataReadRequest_bits_outputTag_id,
  input         io_dataWriteRequest_ready,
  output        io_dataWriteRequest_valid,
  output [63:0] io_dataWriteRequest_bits_address,
  output [63:0] io_dataWriteRequest_bits_data,
  output [7:0]  io_dataWriteRequest_bits_mask
);
  wire  inputArbiter_clock; // @[DataMemoryBuffer.scala 28:36]
  wire  inputArbiter_reset; // @[DataMemoryBuffer.scala 28:36]
  wire  inputArbiter_io_in_0_ready; // @[DataMemoryBuffer.scala 28:36]
  wire  inputArbiter_io_in_0_valid; // @[DataMemoryBuffer.scala 28:36]
  wire [63:0] inputArbiter_io_in_0_bits_address; // @[DataMemoryBuffer.scala 28:36]
  wire  inputArbiter_io_in_0_bits_tag_threadId; // @[DataMemoryBuffer.scala 28:36]
  wire [3:0] inputArbiter_io_in_0_bits_tag_id; // @[DataMemoryBuffer.scala 28:36]
  wire [63:0] inputArbiter_io_in_0_bits_data; // @[DataMemoryBuffer.scala 28:36]
  wire  inputArbiter_io_in_0_bits_accessInfo_accessType; // @[DataMemoryBuffer.scala 28:36]
  wire  inputArbiter_io_in_0_bits_accessInfo_signed; // @[DataMemoryBuffer.scala 28:36]
  wire [1:0] inputArbiter_io_in_0_bits_accessInfo_accessWidth; // @[DataMemoryBuffer.scala 28:36]
  wire  inputArbiter_io_in_1_ready; // @[DataMemoryBuffer.scala 28:36]
  wire  inputArbiter_io_in_1_valid; // @[DataMemoryBuffer.scala 28:36]
  wire [63:0] inputArbiter_io_in_1_bits_address; // @[DataMemoryBuffer.scala 28:36]
  wire  inputArbiter_io_in_1_bits_tag_threadId; // @[DataMemoryBuffer.scala 28:36]
  wire [3:0] inputArbiter_io_in_1_bits_tag_id; // @[DataMemoryBuffer.scala 28:36]
  wire [63:0] inputArbiter_io_in_1_bits_data; // @[DataMemoryBuffer.scala 28:36]
  wire  inputArbiter_io_in_1_bits_accessInfo_accessType; // @[DataMemoryBuffer.scala 28:36]
  wire  inputArbiter_io_in_1_bits_accessInfo_signed; // @[DataMemoryBuffer.scala 28:36]
  wire [1:0] inputArbiter_io_in_1_bits_accessInfo_accessWidth; // @[DataMemoryBuffer.scala 28:36]
  wire  inputArbiter_io_out_ready; // @[DataMemoryBuffer.scala 28:36]
  wire  inputArbiter_io_out_valid; // @[DataMemoryBuffer.scala 28:36]
  wire [63:0] inputArbiter_io_out_bits_address; // @[DataMemoryBuffer.scala 28:36]
  wire  inputArbiter_io_out_bits_tag_threadId; // @[DataMemoryBuffer.scala 28:36]
  wire [3:0] inputArbiter_io_out_bits_tag_id; // @[DataMemoryBuffer.scala 28:36]
  wire [63:0] inputArbiter_io_out_bits_data; // @[DataMemoryBuffer.scala 28:36]
  wire  inputArbiter_io_out_bits_accessInfo_accessType; // @[DataMemoryBuffer.scala 28:36]
  wire  inputArbiter_io_out_bits_accessInfo_signed; // @[DataMemoryBuffer.scala 28:36]
  wire [1:0] inputArbiter_io_out_bits_accessInfo_accessWidth; // @[DataMemoryBuffer.scala 28:36]
  wire  inputArbiter_io_chosen; // @[DataMemoryBuffer.scala 28:36]
  wire  buffer_clock; // @[DataMemoryBuffer.scala 34:30]
  wire  buffer_reset; // @[DataMemoryBuffer.scala 34:30]
  wire  buffer_input_ready; // @[DataMemoryBuffer.scala 34:30]
  wire  buffer_input_valid; // @[DataMemoryBuffer.scala 34:30]
  wire [63:0] buffer_input_bits_address; // @[DataMemoryBuffer.scala 34:30]
  wire  buffer_input_bits_tag_threadId; // @[DataMemoryBuffer.scala 34:30]
  wire [3:0] buffer_input_bits_tag_id; // @[DataMemoryBuffer.scala 34:30]
  wire [63:0] buffer_input_bits_data; // @[DataMemoryBuffer.scala 34:30]
  wire  buffer_input_bits_accessInfo_accessType; // @[DataMemoryBuffer.scala 34:30]
  wire  buffer_input_bits_accessInfo_signed; // @[DataMemoryBuffer.scala 34:30]
  wire [1:0] buffer_input_bits_accessInfo_accessWidth; // @[DataMemoryBuffer.scala 34:30]
  wire  buffer_output_ready; // @[DataMemoryBuffer.scala 34:30]
  wire [63:0] buffer_output_bits_address; // @[DataMemoryBuffer.scala 34:30]
  wire  buffer_output_bits_tag_threadId; // @[DataMemoryBuffer.scala 34:30]
  wire [3:0] buffer_output_bits_tag_id; // @[DataMemoryBuffer.scala 34:30]
  wire [63:0] buffer_output_bits_data; // @[DataMemoryBuffer.scala 34:30]
  wire  buffer_output_bits_accessInfo_accessType; // @[DataMemoryBuffer.scala 34:30]
  wire  buffer_output_bits_accessInfo_signed; // @[DataMemoryBuffer.scala 34:30]
  wire [1:0] buffer_output_bits_accessInfo_accessWidth; // @[DataMemoryBuffer.scala 34:30]
  wire  buffer_empty; // @[DataMemoryBuffer.scala 34:30]
  wire  _T_1 = buffer_output_bits_accessInfo_accessType; // @[DataMemoryBuffer.scala 48:38]
  wire  _T_2 = ~buffer_output_bits_accessInfo_accessType; // @[DataMemoryBuffer.scala 57:44]
  wire [60:0] addressUpper = buffer_output_bits_address[63:3]; // @[DataMemoryBuffer.scala 59:39]
  wire [2:0] addressLower = buffer_output_bits_address[2:0]; // @[DataMemoryBuffer.scala 60:39]
  wire [1:0] _io_dataWriteRequest_bits_data_T = buffer_output_bits_accessInfo_accessWidth; // @[DataMemoryBuffer.scala 64:38]
  wire  _io_dataWriteRequest_bits_data_T_2 = addressLower == 3'h0; // @[DataMemoryBuffer.scala 69:29]
  wire  _io_dataWriteRequest_bits_data_T_5 = addressLower == 3'h1; // @[DataMemoryBuffer.scala 69:29]
  wire [15:0] _io_dataWriteRequest_bits_data_T_7 = {buffer_output_bits_data[7:0], 8'h0}; // @[DataMemoryBuffer.scala 69:59]
  wire  _io_dataWriteRequest_bits_data_T_8 = addressLower == 3'h2; // @[DataMemoryBuffer.scala 69:29]
  wire [23:0] _io_dataWriteRequest_bits_data_T_10 = {buffer_output_bits_data[7:0], 16'h0}; // @[DataMemoryBuffer.scala 69:59]
  wire  _io_dataWriteRequest_bits_data_T_11 = addressLower == 3'h3; // @[DataMemoryBuffer.scala 69:29]
  wire [31:0] _io_dataWriteRequest_bits_data_T_13 = {buffer_output_bits_data[7:0], 24'h0}; // @[DataMemoryBuffer.scala 69:59]
  wire  _io_dataWriteRequest_bits_data_T_14 = addressLower == 3'h4; // @[DataMemoryBuffer.scala 69:29]
  wire [39:0] _io_dataWriteRequest_bits_data_T_16 = {buffer_output_bits_data[7:0], 32'h0}; // @[DataMemoryBuffer.scala 69:59]
  wire  _io_dataWriteRequest_bits_data_T_17 = addressLower == 3'h5; // @[DataMemoryBuffer.scala 69:29]
  wire [47:0] _io_dataWriteRequest_bits_data_T_19 = {buffer_output_bits_data[7:0], 40'h0}; // @[DataMemoryBuffer.scala 69:59]
  wire  _io_dataWriteRequest_bits_data_T_20 = addressLower == 3'h6; // @[DataMemoryBuffer.scala 69:29]
  wire [55:0] _io_dataWriteRequest_bits_data_T_22 = {buffer_output_bits_data[7:0], 48'h0}; // @[DataMemoryBuffer.scala 69:59]
  wire  _io_dataWriteRequest_bits_data_T_23 = addressLower == 3'h7; // @[DataMemoryBuffer.scala 69:29]
  wire [63:0] _io_dataWriteRequest_bits_data_T_25 = {buffer_output_bits_data[7:0], 56'h0}; // @[DataMemoryBuffer.scala 69:59]
  wire [7:0] _io_dataWriteRequest_bits_data_T_26 = _io_dataWriteRequest_bits_data_T_2 ? buffer_output_bits_data[7:0] : 8'h0
    ; // @[Mux.scala 27:73]
  wire [15:0] _io_dataWriteRequest_bits_data_T_27 = _io_dataWriteRequest_bits_data_T_5 ?
    _io_dataWriteRequest_bits_data_T_7 : 16'h0; // @[Mux.scala 27:73]
  wire [23:0] _io_dataWriteRequest_bits_data_T_28 = _io_dataWriteRequest_bits_data_T_8 ?
    _io_dataWriteRequest_bits_data_T_10 : 24'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_dataWriteRequest_bits_data_T_29 = _io_dataWriteRequest_bits_data_T_11 ?
    _io_dataWriteRequest_bits_data_T_13 : 32'h0; // @[Mux.scala 27:73]
  wire [39:0] _io_dataWriteRequest_bits_data_T_30 = _io_dataWriteRequest_bits_data_T_14 ?
    _io_dataWriteRequest_bits_data_T_16 : 40'h0; // @[Mux.scala 27:73]
  wire [47:0] _io_dataWriteRequest_bits_data_T_31 = _io_dataWriteRequest_bits_data_T_17 ?
    _io_dataWriteRequest_bits_data_T_19 : 48'h0; // @[Mux.scala 27:73]
  wire [55:0] _io_dataWriteRequest_bits_data_T_32 = _io_dataWriteRequest_bits_data_T_20 ?
    _io_dataWriteRequest_bits_data_T_22 : 56'h0; // @[Mux.scala 27:73]
  wire [63:0] _io_dataWriteRequest_bits_data_T_33 = _io_dataWriteRequest_bits_data_T_23 ?
    _io_dataWriteRequest_bits_data_T_25 : 64'h0; // @[Mux.scala 27:73]
  wire [15:0] _GEN_35 = {{8'd0}, _io_dataWriteRequest_bits_data_T_26}; // @[Mux.scala 27:73]
  wire [15:0] _io_dataWriteRequest_bits_data_T_34 = _GEN_35 | _io_dataWriteRequest_bits_data_T_27; // @[Mux.scala 27:73]
  wire [23:0] _GEN_36 = {{8'd0}, _io_dataWriteRequest_bits_data_T_34}; // @[Mux.scala 27:73]
  wire [23:0] _io_dataWriteRequest_bits_data_T_35 = _GEN_36 | _io_dataWriteRequest_bits_data_T_28; // @[Mux.scala 27:73]
  wire [31:0] _GEN_37 = {{8'd0}, _io_dataWriteRequest_bits_data_T_35}; // @[Mux.scala 27:73]
  wire [31:0] _io_dataWriteRequest_bits_data_T_36 = _GEN_37 | _io_dataWriteRequest_bits_data_T_29; // @[Mux.scala 27:73]
  wire [39:0] _GEN_38 = {{8'd0}, _io_dataWriteRequest_bits_data_T_36}; // @[Mux.scala 27:73]
  wire [39:0] _io_dataWriteRequest_bits_data_T_37 = _GEN_38 | _io_dataWriteRequest_bits_data_T_30; // @[Mux.scala 27:73]
  wire [47:0] _GEN_39 = {{8'd0}, _io_dataWriteRequest_bits_data_T_37}; // @[Mux.scala 27:73]
  wire [47:0] _io_dataWriteRequest_bits_data_T_38 = _GEN_39 | _io_dataWriteRequest_bits_data_T_31; // @[Mux.scala 27:73]
  wire [55:0] _GEN_40 = {{8'd0}, _io_dataWriteRequest_bits_data_T_38}; // @[Mux.scala 27:73]
  wire [55:0] _io_dataWriteRequest_bits_data_T_39 = _GEN_40 | _io_dataWriteRequest_bits_data_T_32; // @[Mux.scala 27:73]
  wire [63:0] _GEN_41 = {{8'd0}, _io_dataWriteRequest_bits_data_T_39}; // @[Mux.scala 27:73]
  wire [63:0] _io_dataWriteRequest_bits_data_T_40 = _GEN_41 | _io_dataWriteRequest_bits_data_T_33; // @[Mux.scala 27:73]
  wire  _io_dataWriteRequest_bits_data_T_43 = addressLower[2:1] == 2'h0; // @[DataMemoryBuffer.scala 74:35]
  wire  _io_dataWriteRequest_bits_data_T_47 = addressLower[2:1] == 2'h1; // @[DataMemoryBuffer.scala 74:35]
  wire [31:0] _io_dataWriteRequest_bits_data_T_49 = {buffer_output_bits_data[15:0], 16'h0}; // @[DataMemoryBuffer.scala 74:66]
  wire  _io_dataWriteRequest_bits_data_T_51 = addressLower[2:1] == 2'h2; // @[DataMemoryBuffer.scala 74:35]
  wire [47:0] _io_dataWriteRequest_bits_data_T_53 = {buffer_output_bits_data[15:0], 32'h0}; // @[DataMemoryBuffer.scala 74:66]
  wire  _io_dataWriteRequest_bits_data_T_55 = addressLower[2:1] == 2'h3; // @[DataMemoryBuffer.scala 74:35]
  wire [63:0] _io_dataWriteRequest_bits_data_T_57 = {buffer_output_bits_data[15:0], 48'h0}; // @[DataMemoryBuffer.scala 74:66]
  wire [15:0] _io_dataWriteRequest_bits_data_T_58 = _io_dataWriteRequest_bits_data_T_43 ? buffer_output_bits_data[15:0]
     : 16'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_dataWriteRequest_bits_data_T_59 = _io_dataWriteRequest_bits_data_T_47 ?
    _io_dataWriteRequest_bits_data_T_49 : 32'h0; // @[Mux.scala 27:73]
  wire [47:0] _io_dataWriteRequest_bits_data_T_60 = _io_dataWriteRequest_bits_data_T_51 ?
    _io_dataWriteRequest_bits_data_T_53 : 48'h0; // @[Mux.scala 27:73]
  wire [63:0] _io_dataWriteRequest_bits_data_T_61 = _io_dataWriteRequest_bits_data_T_55 ?
    _io_dataWriteRequest_bits_data_T_57 : 64'h0; // @[Mux.scala 27:73]
  wire [31:0] _GEN_42 = {{16'd0}, _io_dataWriteRequest_bits_data_T_58}; // @[Mux.scala 27:73]
  wire [31:0] _io_dataWriteRequest_bits_data_T_62 = _GEN_42 | _io_dataWriteRequest_bits_data_T_59; // @[Mux.scala 27:73]
  wire [47:0] _GEN_43 = {{16'd0}, _io_dataWriteRequest_bits_data_T_62}; // @[Mux.scala 27:73]
  wire [47:0] _io_dataWriteRequest_bits_data_T_63 = _GEN_43 | _io_dataWriteRequest_bits_data_T_60; // @[Mux.scala 27:73]
  wire [63:0] _GEN_44 = {{16'd0}, _io_dataWriteRequest_bits_data_T_63}; // @[Mux.scala 27:73]
  wire [63:0] _io_dataWriteRequest_bits_data_T_64 = _GEN_44 | _io_dataWriteRequest_bits_data_T_61; // @[Mux.scala 27:73]
  wire  _io_dataWriteRequest_bits_data_T_67 = ~addressLower[2]; // @[DataMemoryBuffer.scala 79:32]
  wire [63:0] _io_dataWriteRequest_bits_data_T_73 = {buffer_output_bits_data[31:0], 32'h0}; // @[DataMemoryBuffer.scala 79:63]
  wire [31:0] _io_dataWriteRequest_bits_data_T_74 = _io_dataWriteRequest_bits_data_T_67 ? buffer_output_bits_data[31:0]
     : 32'h0; // @[Mux.scala 27:73]
  wire [63:0] _io_dataWriteRequest_bits_data_T_75 = addressLower[2] ? _io_dataWriteRequest_bits_data_T_73 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _GEN_45 = {{32'd0}, _io_dataWriteRequest_bits_data_T_74}; // @[Mux.scala 27:73]
  wire [63:0] _io_dataWriteRequest_bits_data_T_76 = _GEN_45 | _io_dataWriteRequest_bits_data_T_75; // @[Mux.scala 27:73]
  wire [63:0] _io_dataWriteRequest_bits_data_T_79 = 2'h0 == _io_dataWriteRequest_bits_data_T ?
    _io_dataWriteRequest_bits_data_T_40 : 64'h0; // @[Mux.scala 81:58]
  wire [63:0] _io_dataWriteRequest_bits_data_T_81 = 2'h1 == _io_dataWriteRequest_bits_data_T ?
    _io_dataWriteRequest_bits_data_T_64 : _io_dataWriteRequest_bits_data_T_79; // @[Mux.scala 81:58]
  wire [63:0] _io_dataWriteRequest_bits_data_T_83 = 2'h2 == _io_dataWriteRequest_bits_data_T ?
    _io_dataWriteRequest_bits_data_T_76 : _io_dataWriteRequest_bits_data_T_81; // @[Mux.scala 81:58]
  wire [1:0] _io_dataWriteRequest_bits_mask_T_11 = _io_dataWriteRequest_bits_data_T_5 ? 2'h2 : 2'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_dataWriteRequest_bits_mask_T_12 = _io_dataWriteRequest_bits_data_T_8 ? 3'h4 : 3'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_dataWriteRequest_bits_mask_T_13 = _io_dataWriteRequest_bits_data_T_11 ? 4'h8 : 4'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_dataWriteRequest_bits_mask_T_14 = _io_dataWriteRequest_bits_data_T_14 ? 5'h10 : 5'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_dataWriteRequest_bits_mask_T_15 = _io_dataWriteRequest_bits_data_T_17 ? 6'h20 : 6'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_dataWriteRequest_bits_mask_T_16 = _io_dataWriteRequest_bits_data_T_20 ? 7'h40 : 7'h0; // @[Mux.scala 27:73]
  wire [7:0] _io_dataWriteRequest_bits_mask_T_17 = _io_dataWriteRequest_bits_data_T_23 ? 8'h80 : 8'h0; // @[Mux.scala 27:73]
  wire [1:0] _GEN_46 = {{1'd0}, _io_dataWriteRequest_bits_data_T_2}; // @[Mux.scala 27:73]
  wire [1:0] _io_dataWriteRequest_bits_mask_T_18 = _GEN_46 | _io_dataWriteRequest_bits_mask_T_11; // @[Mux.scala 27:73]
  wire [2:0] _GEN_47 = {{1'd0}, _io_dataWriteRequest_bits_mask_T_18}; // @[Mux.scala 27:73]
  wire [2:0] _io_dataWriteRequest_bits_mask_T_19 = _GEN_47 | _io_dataWriteRequest_bits_mask_T_12; // @[Mux.scala 27:73]
  wire [3:0] _GEN_48 = {{1'd0}, _io_dataWriteRequest_bits_mask_T_19}; // @[Mux.scala 27:73]
  wire [3:0] _io_dataWriteRequest_bits_mask_T_20 = _GEN_48 | _io_dataWriteRequest_bits_mask_T_13; // @[Mux.scala 27:73]
  wire [4:0] _GEN_49 = {{1'd0}, _io_dataWriteRequest_bits_mask_T_20}; // @[Mux.scala 27:73]
  wire [4:0] _io_dataWriteRequest_bits_mask_T_21 = _GEN_49 | _io_dataWriteRequest_bits_mask_T_14; // @[Mux.scala 27:73]
  wire [5:0] _GEN_50 = {{1'd0}, _io_dataWriteRequest_bits_mask_T_21}; // @[Mux.scala 27:73]
  wire [5:0] _io_dataWriteRequest_bits_mask_T_22 = _GEN_50 | _io_dataWriteRequest_bits_mask_T_15; // @[Mux.scala 27:73]
  wire [6:0] _GEN_51 = {{1'd0}, _io_dataWriteRequest_bits_mask_T_22}; // @[Mux.scala 27:73]
  wire [6:0] _io_dataWriteRequest_bits_mask_T_23 = _GEN_51 | _io_dataWriteRequest_bits_mask_T_16; // @[Mux.scala 27:73]
  wire [7:0] _GEN_52 = {{1'd0}, _io_dataWriteRequest_bits_mask_T_23}; // @[Mux.scala 27:73]
  wire [7:0] _io_dataWriteRequest_bits_mask_T_24 = _GEN_52 | _io_dataWriteRequest_bits_mask_T_17; // @[Mux.scala 27:73]
  wire [1:0] _io_dataWriteRequest_bits_mask_T_34 = _io_dataWriteRequest_bits_data_T_43 ? 2'h3 : 2'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_dataWriteRequest_bits_mask_T_35 = _io_dataWriteRequest_bits_data_T_47 ? 4'hc : 4'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_dataWriteRequest_bits_mask_T_36 = _io_dataWriteRequest_bits_data_T_51 ? 6'h30 : 6'h0; // @[Mux.scala 27:73]
  wire [7:0] _io_dataWriteRequest_bits_mask_T_37 = _io_dataWriteRequest_bits_data_T_55 ? 8'hc0 : 8'h0; // @[Mux.scala 27:73]
  wire [3:0] _GEN_53 = {{2'd0}, _io_dataWriteRequest_bits_mask_T_34}; // @[Mux.scala 27:73]
  wire [3:0] _io_dataWriteRequest_bits_mask_T_38 = _GEN_53 | _io_dataWriteRequest_bits_mask_T_35; // @[Mux.scala 27:73]
  wire [5:0] _GEN_54 = {{2'd0}, _io_dataWriteRequest_bits_mask_T_38}; // @[Mux.scala 27:73]
  wire [5:0] _io_dataWriteRequest_bits_mask_T_39 = _GEN_54 | _io_dataWriteRequest_bits_mask_T_36; // @[Mux.scala 27:73]
  wire [7:0] _GEN_55 = {{2'd0}, _io_dataWriteRequest_bits_mask_T_39}; // @[Mux.scala 27:73]
  wire [7:0] _io_dataWriteRequest_bits_mask_T_40 = _GEN_55 | _io_dataWriteRequest_bits_mask_T_37; // @[Mux.scala 27:73]
  wire [3:0] _io_dataWriteRequest_bits_mask_T_46 = _io_dataWriteRequest_bits_data_T_67 ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [7:0] _io_dataWriteRequest_bits_mask_T_47 = addressLower[2] ? 8'hf0 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _GEN_56 = {{4'd0}, _io_dataWriteRequest_bits_mask_T_46}; // @[Mux.scala 27:73]
  wire [7:0] _io_dataWriteRequest_bits_mask_T_48 = _GEN_56 | _io_dataWriteRequest_bits_mask_T_47; // @[Mux.scala 27:73]
  wire [7:0] _io_dataWriteRequest_bits_mask_T_51 = 2'h0 == _io_dataWriteRequest_bits_data_T ?
    _io_dataWriteRequest_bits_mask_T_24 : 8'h0; // @[Mux.scala 81:58]
  wire [7:0] _io_dataWriteRequest_bits_mask_T_53 = 2'h1 == _io_dataWriteRequest_bits_data_T ?
    _io_dataWriteRequest_bits_mask_T_40 : _io_dataWriteRequest_bits_mask_T_51; // @[Mux.scala 81:58]
  wire [7:0] _io_dataWriteRequest_bits_mask_T_55 = 2'h2 == _io_dataWriteRequest_bits_data_T ?
    _io_dataWriteRequest_bits_mask_T_48 : _io_dataWriteRequest_bits_mask_T_53; // @[Mux.scala 81:58]
  wire  _GEN_4 = buffer_output_bits_tag_threadId; // @[DataMemoryBuffer.scala 57:72 62:42]
  wire [3:0] _GEN_5 = buffer_output_bits_tag_id; // @[DataMemoryBuffer.scala 57:72 62:42]
  wire  _GEN_8 = ~buffer_output_bits_accessInfo_accessType & io_dataWriteRequest_ready; // @[DataMemoryBuffer.scala 38:23 57:72]
  wire  _GEN_15 = buffer_output_bits_accessInfo_accessType ? io_dataReadRequest_ready : _GEN_8; // @[DataMemoryBuffer.scala 48:65]
  wire  _GEN_16 = buffer_output_bits_accessInfo_accessType ? 1'h0 : _T_2; // @[DataMemoryBuffer.scala 44:29 48:65]
  B4RRArbiter inputArbiter ( // @[DataMemoryBuffer.scala 28:36]
    .clock(inputArbiter_clock),
    .reset(inputArbiter_reset),
    .io_in_0_ready(inputArbiter_io_in_0_ready),
    .io_in_0_valid(inputArbiter_io_in_0_valid),
    .io_in_0_bits_address(inputArbiter_io_in_0_bits_address),
    .io_in_0_bits_tag_threadId(inputArbiter_io_in_0_bits_tag_threadId),
    .io_in_0_bits_tag_id(inputArbiter_io_in_0_bits_tag_id),
    .io_in_0_bits_data(inputArbiter_io_in_0_bits_data),
    .io_in_0_bits_accessInfo_accessType(inputArbiter_io_in_0_bits_accessInfo_accessType),
    .io_in_0_bits_accessInfo_signed(inputArbiter_io_in_0_bits_accessInfo_signed),
    .io_in_0_bits_accessInfo_accessWidth(inputArbiter_io_in_0_bits_accessInfo_accessWidth),
    .io_in_1_ready(inputArbiter_io_in_1_ready),
    .io_in_1_valid(inputArbiter_io_in_1_valid),
    .io_in_1_bits_address(inputArbiter_io_in_1_bits_address),
    .io_in_1_bits_tag_threadId(inputArbiter_io_in_1_bits_tag_threadId),
    .io_in_1_bits_tag_id(inputArbiter_io_in_1_bits_tag_id),
    .io_in_1_bits_data(inputArbiter_io_in_1_bits_data),
    .io_in_1_bits_accessInfo_accessType(inputArbiter_io_in_1_bits_accessInfo_accessType),
    .io_in_1_bits_accessInfo_signed(inputArbiter_io_in_1_bits_accessInfo_signed),
    .io_in_1_bits_accessInfo_accessWidth(inputArbiter_io_in_1_bits_accessInfo_accessWidth),
    .io_out_ready(inputArbiter_io_out_ready),
    .io_out_valid(inputArbiter_io_out_valid),
    .io_out_bits_address(inputArbiter_io_out_bits_address),
    .io_out_bits_tag_threadId(inputArbiter_io_out_bits_tag_threadId),
    .io_out_bits_tag_id(inputArbiter_io_out_bits_tag_id),
    .io_out_bits_data(inputArbiter_io_out_bits_data),
    .io_out_bits_accessInfo_accessType(inputArbiter_io_out_bits_accessInfo_accessType),
    .io_out_bits_accessInfo_signed(inputArbiter_io_out_bits_accessInfo_signed),
    .io_out_bits_accessInfo_accessWidth(inputArbiter_io_out_bits_accessInfo_accessWidth),
    .io_chosen(inputArbiter_io_chosen)
  );
  FIFO buffer ( // @[DataMemoryBuffer.scala 34:30]
    .clock(buffer_clock),
    .reset(buffer_reset),
    .input_ready(buffer_input_ready),
    .input_valid(buffer_input_valid),
    .input_bits_address(buffer_input_bits_address),
    .input_bits_tag_threadId(buffer_input_bits_tag_threadId),
    .input_bits_tag_id(buffer_input_bits_tag_id),
    .input_bits_data(buffer_input_bits_data),
    .input_bits_accessInfo_accessType(buffer_input_bits_accessInfo_accessType),
    .input_bits_accessInfo_signed(buffer_input_bits_accessInfo_signed),
    .input_bits_accessInfo_accessWidth(buffer_input_bits_accessInfo_accessWidth),
    .output_ready(buffer_output_ready),
    .output_bits_address(buffer_output_bits_address),
    .output_bits_tag_threadId(buffer_output_bits_tag_threadId),
    .output_bits_tag_id(buffer_output_bits_tag_id),
    .output_bits_data(buffer_output_bits_data),
    .output_bits_accessInfo_accessType(buffer_output_bits_accessInfo_accessType),
    .output_bits_accessInfo_signed(buffer_output_bits_accessInfo_signed),
    .output_bits_accessInfo_accessWidth(buffer_output_bits_accessInfo_accessWidth),
    .empty(buffer_empty)
  );
  assign io_dataIn_0_ready = inputArbiter_io_in_0_ready; // @[DataMemoryBuffer.scala 32:29]
  assign io_dataIn_1_ready = inputArbiter_io_in_1_ready; // @[DataMemoryBuffer.scala 32:29]
  assign io_dataReadRequest_valid = ~buffer_empty & _T_1; // @[DataMemoryBuffer.scala 46:23 42:28]
  assign io_dataReadRequest_bits_address = buffer_output_bits_address; // @[DataMemoryBuffer.scala 48:65 50:39]
  assign io_dataReadRequest_bits_size = buffer_output_bits_accessInfo_accessWidth; // @[DataMemoryBuffer.scala 48:65 51:36]
  assign io_dataReadRequest_bits_signed = buffer_output_bits_accessInfo_signed; // @[DataMemoryBuffer.scala 48:65 53:38]
  assign io_dataReadRequest_bits_outputTag_threadId = buffer_output_bits_accessInfo_accessType ?
    buffer_output_bits_tag_threadId : _GEN_4; // @[DataMemoryBuffer.scala 48:65 52:41]
  assign io_dataReadRequest_bits_outputTag_id = buffer_output_bits_accessInfo_accessType ? buffer_output_bits_tag_id :
    _GEN_5; // @[DataMemoryBuffer.scala 48:65 52:41]
  assign io_dataWriteRequest_valid = ~buffer_empty & _GEN_16; // @[DataMemoryBuffer.scala 46:23 44:29]
  assign io_dataWriteRequest_bits_address = {addressUpper,3'h0}; // @[DataMemoryBuffer.scala 61:56]
  assign io_dataWriteRequest_bits_data = 2'h3 == _io_dataWriteRequest_bits_data_T ? buffer_output_bits_data :
    _io_dataWriteRequest_bits_data_T_83; // @[Mux.scala 81:58]
  assign io_dataWriteRequest_bits_mask = 2'h3 == _io_dataWriteRequest_bits_data_T ? 8'hff :
    _io_dataWriteRequest_bits_mask_T_55; // @[Mux.scala 81:58]
  assign inputArbiter_clock = clock;
  assign inputArbiter_reset = reset;
  assign inputArbiter_io_in_0_valid = io_dataIn_0_valid; // @[DataMemoryBuffer.scala 32:29]
  assign inputArbiter_io_in_0_bits_address = io_dataIn_0_bits_address; // @[DataMemoryBuffer.scala 32:29]
  assign inputArbiter_io_in_0_bits_tag_threadId = io_dataIn_0_bits_tag_threadId; // @[DataMemoryBuffer.scala 32:29]
  assign inputArbiter_io_in_0_bits_tag_id = io_dataIn_0_bits_tag_id; // @[DataMemoryBuffer.scala 32:29]
  assign inputArbiter_io_in_0_bits_data = io_dataIn_0_bits_data; // @[DataMemoryBuffer.scala 32:29]
  assign inputArbiter_io_in_0_bits_accessInfo_accessType = io_dataIn_0_bits_accessInfo_accessType; // @[DataMemoryBuffer.scala 32:29]
  assign inputArbiter_io_in_0_bits_accessInfo_signed = io_dataIn_0_bits_accessInfo_signed; // @[DataMemoryBuffer.scala 32:29]
  assign inputArbiter_io_in_0_bits_accessInfo_accessWidth = io_dataIn_0_bits_accessInfo_accessWidth; // @[DataMemoryBuffer.scala 32:29]
  assign inputArbiter_io_in_1_valid = io_dataIn_1_valid; // @[DataMemoryBuffer.scala 32:29]
  assign inputArbiter_io_in_1_bits_address = io_dataIn_1_bits_address; // @[DataMemoryBuffer.scala 32:29]
  assign inputArbiter_io_in_1_bits_tag_threadId = io_dataIn_1_bits_tag_threadId; // @[DataMemoryBuffer.scala 32:29]
  assign inputArbiter_io_in_1_bits_tag_id = io_dataIn_1_bits_tag_id; // @[DataMemoryBuffer.scala 32:29]
  assign inputArbiter_io_in_1_bits_data = io_dataIn_1_bits_data; // @[DataMemoryBuffer.scala 32:29]
  assign inputArbiter_io_in_1_bits_accessInfo_accessType = io_dataIn_1_bits_accessInfo_accessType; // @[DataMemoryBuffer.scala 32:29]
  assign inputArbiter_io_in_1_bits_accessInfo_signed = io_dataIn_1_bits_accessInfo_signed; // @[DataMemoryBuffer.scala 32:29]
  assign inputArbiter_io_in_1_bits_accessInfo_accessWidth = io_dataIn_1_bits_accessInfo_accessWidth; // @[DataMemoryBuffer.scala 32:29]
  assign inputArbiter_io_out_ready = buffer_input_ready; // @[DataMemoryBuffer.scala 37:16]
  assign buffer_clock = clock;
  assign buffer_reset = reset;
  assign buffer_input_valid = inputArbiter_io_out_valid; // @[DataMemoryBuffer.scala 37:16]
  assign buffer_input_bits_address = inputArbiter_io_out_bits_address; // @[DataMemoryBuffer.scala 37:16]
  assign buffer_input_bits_tag_threadId = inputArbiter_io_out_bits_tag_threadId; // @[DataMemoryBuffer.scala 37:16]
  assign buffer_input_bits_tag_id = inputArbiter_io_out_bits_tag_id; // @[DataMemoryBuffer.scala 37:16]
  assign buffer_input_bits_data = inputArbiter_io_out_bits_data; // @[DataMemoryBuffer.scala 37:16]
  assign buffer_input_bits_accessInfo_accessType = inputArbiter_io_out_bits_accessInfo_accessType; // @[DataMemoryBuffer.scala 37:16]
  assign buffer_input_bits_accessInfo_signed = inputArbiter_io_out_bits_accessInfo_signed; // @[DataMemoryBuffer.scala 37:16]
  assign buffer_input_bits_accessInfo_accessWidth = inputArbiter_io_out_bits_accessInfo_accessWidth; // @[DataMemoryBuffer.scala 37:16]
  assign buffer_output_ready = ~buffer_empty & _GEN_15; // @[DataMemoryBuffer.scala 38:23 46:23]
endmodule
module Queue_1(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input         io_enq_bits_resultType,
  input  [63:0] io_enq_bits_value,
  input         io_enq_bits_isError,
  input         io_enq_bits_tag_threadId,
  input  [3:0]  io_enq_bits_tag_id,
  output        io_deq_valid,
  output        io_deq_bits_resultType,
  output [63:0] io_deq_bits_value,
  output        io_deq_bits_isError,
  output        io_deq_bits_tag_threadId,
  output [3:0]  io_deq_bits_tag_id,
  input         io_flush
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_12;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
`endif // RANDOMIZE_REG_INIT
  reg  ram_resultType [0:7]; // @[Decoupled.scala 273:44]
  wire  ram_resultType_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:44]
  wire [2:0] ram_resultType_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:44]
  wire  ram_resultType_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:44]
  wire  ram_resultType_MPORT_data; // @[Decoupled.scala 273:44]
  wire [2:0] ram_resultType_MPORT_addr; // @[Decoupled.scala 273:44]
  wire  ram_resultType_MPORT_mask; // @[Decoupled.scala 273:44]
  wire  ram_resultType_MPORT_en; // @[Decoupled.scala 273:44]
  reg  ram_resultType_io_deq_bits_MPORT_en_pipe_0;
  reg [2:0] ram_resultType_io_deq_bits_MPORT_addr_pipe_0;
  reg [63:0] ram_value [0:7]; // @[Decoupled.scala 273:44]
  wire  ram_value_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:44]
  wire [2:0] ram_value_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:44]
  wire [63:0] ram_value_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:44]
  wire [63:0] ram_value_MPORT_data; // @[Decoupled.scala 273:44]
  wire [2:0] ram_value_MPORT_addr; // @[Decoupled.scala 273:44]
  wire  ram_value_MPORT_mask; // @[Decoupled.scala 273:44]
  wire  ram_value_MPORT_en; // @[Decoupled.scala 273:44]
  reg  ram_value_io_deq_bits_MPORT_en_pipe_0;
  reg [2:0] ram_value_io_deq_bits_MPORT_addr_pipe_0;
  reg  ram_isError [0:7]; // @[Decoupled.scala 273:44]
  wire  ram_isError_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:44]
  wire [2:0] ram_isError_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:44]
  wire  ram_isError_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:44]
  wire  ram_isError_MPORT_data; // @[Decoupled.scala 273:44]
  wire [2:0] ram_isError_MPORT_addr; // @[Decoupled.scala 273:44]
  wire  ram_isError_MPORT_mask; // @[Decoupled.scala 273:44]
  wire  ram_isError_MPORT_en; // @[Decoupled.scala 273:44]
  reg  ram_isError_io_deq_bits_MPORT_en_pipe_0;
  reg [2:0] ram_isError_io_deq_bits_MPORT_addr_pipe_0;
  reg  ram_tag_threadId [0:7]; // @[Decoupled.scala 273:44]
  wire  ram_tag_threadId_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:44]
  wire [2:0] ram_tag_threadId_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:44]
  wire  ram_tag_threadId_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:44]
  wire  ram_tag_threadId_MPORT_data; // @[Decoupled.scala 273:44]
  wire [2:0] ram_tag_threadId_MPORT_addr; // @[Decoupled.scala 273:44]
  wire  ram_tag_threadId_MPORT_mask; // @[Decoupled.scala 273:44]
  wire  ram_tag_threadId_MPORT_en; // @[Decoupled.scala 273:44]
  reg  ram_tag_threadId_io_deq_bits_MPORT_en_pipe_0;
  reg [2:0] ram_tag_threadId_io_deq_bits_MPORT_addr_pipe_0;
  reg [3:0] ram_tag_id [0:7]; // @[Decoupled.scala 273:44]
  wire  ram_tag_id_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:44]
  wire [2:0] ram_tag_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:44]
  wire [3:0] ram_tag_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:44]
  wire [3:0] ram_tag_id_MPORT_data; // @[Decoupled.scala 273:44]
  wire [2:0] ram_tag_id_MPORT_addr; // @[Decoupled.scala 273:44]
  wire  ram_tag_id_MPORT_mask; // @[Decoupled.scala 273:44]
  wire  ram_tag_id_MPORT_en; // @[Decoupled.scala 273:44]
  reg  ram_tag_id_io_deq_bits_MPORT_en_pipe_0;
  reg [2:0] ram_tag_id_io_deq_bits_MPORT_addr_pipe_0;
  reg [2:0] enq_ptr_value; // @[Counter.scala 61:40]
  reg [2:0] deq_ptr_value; // @[Counter.scala 61:40]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 277:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 278:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 279:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _value_T_1 = enq_ptr_value + 3'h1; // @[Counter.scala 77:24]
  wire [2:0] _value_T_3 = deq_ptr_value + 3'h1; // @[Counter.scala 77:24]
  wire [3:0] _deq_ptr_next_T_1 = 4'h8 - 4'h1; // @[Decoupled.scala 306:57]
  wire [3:0] _GEN_19 = {{1'd0}, deq_ptr_value}; // @[Decoupled.scala 306:42]
  assign ram_resultType_io_deq_bits_MPORT_en = ram_resultType_io_deq_bits_MPORT_en_pipe_0;
  assign ram_resultType_io_deq_bits_MPORT_addr = ram_resultType_io_deq_bits_MPORT_addr_pipe_0;
  assign ram_resultType_io_deq_bits_MPORT_data = ram_resultType[ram_resultType_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:44]
  assign ram_resultType_MPORT_data = io_enq_bits_resultType;
  assign ram_resultType_MPORT_addr = enq_ptr_value;
  assign ram_resultType_MPORT_mask = 1'h1;
  assign ram_resultType_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_value_io_deq_bits_MPORT_en = ram_value_io_deq_bits_MPORT_en_pipe_0;
  assign ram_value_io_deq_bits_MPORT_addr = ram_value_io_deq_bits_MPORT_addr_pipe_0;
  assign ram_value_io_deq_bits_MPORT_data = ram_value[ram_value_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:44]
  assign ram_value_MPORT_data = io_enq_bits_value;
  assign ram_value_MPORT_addr = enq_ptr_value;
  assign ram_value_MPORT_mask = 1'h1;
  assign ram_value_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_isError_io_deq_bits_MPORT_en = ram_isError_io_deq_bits_MPORT_en_pipe_0;
  assign ram_isError_io_deq_bits_MPORT_addr = ram_isError_io_deq_bits_MPORT_addr_pipe_0;
  assign ram_isError_io_deq_bits_MPORT_data = ram_isError[ram_isError_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:44]
  assign ram_isError_MPORT_data = io_enq_bits_isError;
  assign ram_isError_MPORT_addr = enq_ptr_value;
  assign ram_isError_MPORT_mask = 1'h1;
  assign ram_isError_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_tag_threadId_io_deq_bits_MPORT_en = ram_tag_threadId_io_deq_bits_MPORT_en_pipe_0;
  assign ram_tag_threadId_io_deq_bits_MPORT_addr = ram_tag_threadId_io_deq_bits_MPORT_addr_pipe_0;
  assign ram_tag_threadId_io_deq_bits_MPORT_data = ram_tag_threadId[ram_tag_threadId_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:44]
  assign ram_tag_threadId_MPORT_data = io_enq_bits_tag_threadId;
  assign ram_tag_threadId_MPORT_addr = enq_ptr_value;
  assign ram_tag_threadId_MPORT_mask = 1'h1;
  assign ram_tag_threadId_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_tag_id_io_deq_bits_MPORT_en = ram_tag_id_io_deq_bits_MPORT_en_pipe_0;
  assign ram_tag_id_io_deq_bits_MPORT_addr = ram_tag_id_io_deq_bits_MPORT_addr_pipe_0;
  assign ram_tag_id_io_deq_bits_MPORT_data = ram_tag_id[ram_tag_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:44]
  assign ram_tag_id_MPORT_data = io_enq_bits_tag_id;
  assign ram_tag_id_MPORT_addr = enq_ptr_value;
  assign ram_tag_id_MPORT_mask = 1'h1;
  assign ram_tag_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 303:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 302:19]
  assign io_deq_bits_resultType = ram_resultType_io_deq_bits_MPORT_data; // @[Decoupled.scala 308:17]
  assign io_deq_bits_value = ram_value_io_deq_bits_MPORT_data; // @[Decoupled.scala 308:17]
  assign io_deq_bits_isError = ram_isError_io_deq_bits_MPORT_data; // @[Decoupled.scala 308:17]
  assign io_deq_bits_tag_threadId = ram_tag_threadId_io_deq_bits_MPORT_data; // @[Decoupled.scala 308:17]
  assign io_deq_bits_tag_id = ram_tag_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 308:17]
  always @(posedge clock) begin
    if (ram_resultType_MPORT_en & ram_resultType_MPORT_mask) begin
      ram_resultType[ram_resultType_MPORT_addr] <= ram_resultType_MPORT_data; // @[Decoupled.scala 273:44]
    end
    ram_resultType_io_deq_bits_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (io_deq_valid) begin
        if (_GEN_19 == _deq_ptr_next_T_1) begin // @[Decoupled.scala 306:27]
          ram_resultType_io_deq_bits_MPORT_addr_pipe_0 <= 3'h0;
        end else begin
          ram_resultType_io_deq_bits_MPORT_addr_pipe_0 <= _value_T_3;
        end
      end else begin
        ram_resultType_io_deq_bits_MPORT_addr_pipe_0 <= deq_ptr_value;
      end
    end
    if (ram_value_MPORT_en & ram_value_MPORT_mask) begin
      ram_value[ram_value_MPORT_addr] <= ram_value_MPORT_data; // @[Decoupled.scala 273:44]
    end
    ram_value_io_deq_bits_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (io_deq_valid) begin
        if (_GEN_19 == _deq_ptr_next_T_1) begin // @[Decoupled.scala 306:27]
          ram_value_io_deq_bits_MPORT_addr_pipe_0 <= 3'h0;
        end else begin
          ram_value_io_deq_bits_MPORT_addr_pipe_0 <= _value_T_3;
        end
      end else begin
        ram_value_io_deq_bits_MPORT_addr_pipe_0 <= deq_ptr_value;
      end
    end
    if (ram_isError_MPORT_en & ram_isError_MPORT_mask) begin
      ram_isError[ram_isError_MPORT_addr] <= ram_isError_MPORT_data; // @[Decoupled.scala 273:44]
    end
    ram_isError_io_deq_bits_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (io_deq_valid) begin
        if (_GEN_19 == _deq_ptr_next_T_1) begin // @[Decoupled.scala 306:27]
          ram_isError_io_deq_bits_MPORT_addr_pipe_0 <= 3'h0;
        end else begin
          ram_isError_io_deq_bits_MPORT_addr_pipe_0 <= _value_T_3;
        end
      end else begin
        ram_isError_io_deq_bits_MPORT_addr_pipe_0 <= deq_ptr_value;
      end
    end
    if (ram_tag_threadId_MPORT_en & ram_tag_threadId_MPORT_mask) begin
      ram_tag_threadId[ram_tag_threadId_MPORT_addr] <= ram_tag_threadId_MPORT_data; // @[Decoupled.scala 273:44]
    end
    ram_tag_threadId_io_deq_bits_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (io_deq_valid) begin
        if (_GEN_19 == _deq_ptr_next_T_1) begin // @[Decoupled.scala 306:27]
          ram_tag_threadId_io_deq_bits_MPORT_addr_pipe_0 <= 3'h0;
        end else begin
          ram_tag_threadId_io_deq_bits_MPORT_addr_pipe_0 <= _value_T_3;
        end
      end else begin
        ram_tag_threadId_io_deq_bits_MPORT_addr_pipe_0 <= deq_ptr_value;
      end
    end
    if (ram_tag_id_MPORT_en & ram_tag_id_MPORT_mask) begin
      ram_tag_id[ram_tag_id_MPORT_addr] <= ram_tag_id_MPORT_data; // @[Decoupled.scala 273:44]
    end
    ram_tag_id_io_deq_bits_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (io_deq_valid) begin
        if (_GEN_19 == _deq_ptr_next_T_1) begin // @[Decoupled.scala 306:27]
          ram_tag_id_io_deq_bits_MPORT_addr_pipe_0 <= 3'h0;
        end else begin
          ram_tag_id_io_deq_bits_MPORT_addr_pipe_0 <= _value_T_3;
        end
      end else begin
        ram_tag_id_io_deq_bits_MPORT_addr_pipe_0 <= deq_ptr_value;
      end
    end
    if (reset) begin // @[Counter.scala 61:40]
      enq_ptr_value <= 3'h0; // @[Counter.scala 61:40]
    end else if (io_flush) begin // @[Decoupled.scala 296:15]
      enq_ptr_value <= 3'h0; // @[Counter.scala 98:11]
    end else if (do_enq) begin // @[Decoupled.scala 286:16]
      enq_ptr_value <= _value_T_1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      deq_ptr_value <= 3'h0; // @[Counter.scala 61:40]
    end else if (io_flush) begin // @[Decoupled.scala 296:15]
      deq_ptr_value <= 3'h0; // @[Counter.scala 98:11]
    end else if (io_deq_valid) begin // @[Decoupled.scala 290:16]
      deq_ptr_value <= _value_T_3; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (io_flush) begin // @[Decoupled.scala 296:15]
      maybe_full <= 1'h0; // @[Decoupled.scala 299:16]
    end else if (do_enq != io_deq_valid) begin // @[Decoupled.scala 293:27]
      maybe_full <= do_enq; // @[Decoupled.scala 294:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_resultType[initvar] = _RAND_0[0:0];
  _RAND_3 = {2{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_value[initvar] = _RAND_3[63:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_isError[initvar] = _RAND_6[0:0];
  _RAND_9 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_tag_threadId[initvar] = _RAND_9[0:0];
  _RAND_12 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_tag_id[initvar] = _RAND_12[3:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_resultType_io_deq_bits_MPORT_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  ram_resultType_io_deq_bits_MPORT_addr_pipe_0 = _RAND_2[2:0];
  _RAND_4 = {1{`RANDOM}};
  ram_value_io_deq_bits_MPORT_en_pipe_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  ram_value_io_deq_bits_MPORT_addr_pipe_0 = _RAND_5[2:0];
  _RAND_7 = {1{`RANDOM}};
  ram_isError_io_deq_bits_MPORT_en_pipe_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  ram_isError_io_deq_bits_MPORT_addr_pipe_0 = _RAND_8[2:0];
  _RAND_10 = {1{`RANDOM}};
  ram_tag_threadId_io_deq_bits_MPORT_en_pipe_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  ram_tag_threadId_io_deq_bits_MPORT_addr_pipe_0 = _RAND_11[2:0];
  _RAND_13 = {1{`RANDOM}};
  ram_tag_id_io_deq_bits_MPORT_en_pipe_0 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  ram_tag_id_io_deq_bits_MPORT_addr_pipe_0 = _RAND_14[2:0];
  _RAND_15 = {1{`RANDOM}};
  enq_ptr_value = _RAND_15[2:0];
  _RAND_16 = {1{`RANDOM}};
  deq_ptr_value = _RAND_16[2:0];
  _RAND_17 = {1{`RANDOM}};
  maybe_full = _RAND_17[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module FIFO_1(
  input         clock,
  input         reset,
  output        input_ready,
  input         input_valid,
  input         input_bits_resultType,
  input  [63:0] input_bits_value,
  input         input_bits_isError,
  input         input_bits_tag_threadId,
  input  [3:0]  input_bits_tag_id,
  output        output_valid,
  output        output_bits_resultType,
  output [63:0] output_bits_value,
  output        output_bits_isError,
  output        output_bits_tag_threadId,
  output [3:0]  output_bits_tag_id,
  input         flush
);
  wire  queue_clock; // @[FIFO.scala 16:29]
  wire  queue_reset; // @[FIFO.scala 16:29]
  wire  queue_io_enq_ready; // @[FIFO.scala 16:29]
  wire  queue_io_enq_valid; // @[FIFO.scala 16:29]
  wire  queue_io_enq_bits_resultType; // @[FIFO.scala 16:29]
  wire [63:0] queue_io_enq_bits_value; // @[FIFO.scala 16:29]
  wire  queue_io_enq_bits_isError; // @[FIFO.scala 16:29]
  wire  queue_io_enq_bits_tag_threadId; // @[FIFO.scala 16:29]
  wire [3:0] queue_io_enq_bits_tag_id; // @[FIFO.scala 16:29]
  wire  queue_io_deq_valid; // @[FIFO.scala 16:29]
  wire  queue_io_deq_bits_resultType; // @[FIFO.scala 16:29]
  wire [63:0] queue_io_deq_bits_value; // @[FIFO.scala 16:29]
  wire  queue_io_deq_bits_isError; // @[FIFO.scala 16:29]
  wire  queue_io_deq_bits_tag_threadId; // @[FIFO.scala 16:29]
  wire [3:0] queue_io_deq_bits_tag_id; // @[FIFO.scala 16:29]
  wire  queue_io_flush; // @[FIFO.scala 16:29]
  Queue_1 queue ( // @[FIFO.scala 16:29]
    .clock(queue_clock),
    .reset(queue_reset),
    .io_enq_ready(queue_io_enq_ready),
    .io_enq_valid(queue_io_enq_valid),
    .io_enq_bits_resultType(queue_io_enq_bits_resultType),
    .io_enq_bits_value(queue_io_enq_bits_value),
    .io_enq_bits_isError(queue_io_enq_bits_isError),
    .io_enq_bits_tag_threadId(queue_io_enq_bits_tag_threadId),
    .io_enq_bits_tag_id(queue_io_enq_bits_tag_id),
    .io_deq_valid(queue_io_deq_valid),
    .io_deq_bits_resultType(queue_io_deq_bits_resultType),
    .io_deq_bits_value(queue_io_deq_bits_value),
    .io_deq_bits_isError(queue_io_deq_bits_isError),
    .io_deq_bits_tag_threadId(queue_io_deq_bits_tag_threadId),
    .io_deq_bits_tag_id(queue_io_deq_bits_tag_id),
    .io_flush(queue_io_flush)
  );
  assign input_ready = queue_io_enq_ready; // @[FIFO.scala 19:16]
  assign output_valid = queue_io_deq_valid; // @[FIFO.scala 20:10]
  assign output_bits_resultType = queue_io_deq_bits_resultType; // @[FIFO.scala 20:10]
  assign output_bits_value = queue_io_deq_bits_value; // @[FIFO.scala 20:10]
  assign output_bits_isError = queue_io_deq_bits_isError; // @[FIFO.scala 20:10]
  assign output_bits_tag_threadId = queue_io_deq_bits_tag_threadId; // @[FIFO.scala 20:10]
  assign output_bits_tag_id = queue_io_deq_bits_tag_id; // @[FIFO.scala 20:10]
  assign queue_clock = clock;
  assign queue_reset = reset;
  assign queue_io_enq_valid = input_valid; // @[FIFO.scala 19:16]
  assign queue_io_enq_bits_resultType = input_bits_resultType; // @[FIFO.scala 19:16]
  assign queue_io_enq_bits_value = input_bits_value; // @[FIFO.scala 19:16]
  assign queue_io_enq_bits_isError = input_bits_isError; // @[FIFO.scala 19:16]
  assign queue_io_enq_bits_tag_threadId = input_bits_tag_threadId; // @[FIFO.scala 19:16]
  assign queue_io_enq_bits_tag_id = input_bits_tag_id; // @[FIFO.scala 19:16]
  assign queue_io_flush = flush; // @[FIFO.scala 23:15]
endmodule
module Arbiter(
  output        io_in_0_ready,
  input         io_in_0_valid,
  input         io_in_0_bits_resultType,
  input  [63:0] io_in_0_bits_value,
  input         io_in_0_bits_tag_threadId,
  input  [3:0]  io_in_0_bits_tag_id,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input         io_in_1_bits_resultType,
  input  [63:0] io_in_1_bits_value,
  input         io_in_1_bits_tag_threadId,
  input  [3:0]  io_in_1_bits_tag_id,
  output        io_in_2_ready,
  input         io_in_2_valid,
  input  [63:0] io_in_2_bits_value,
  input         io_in_2_bits_isError,
  input         io_in_2_bits_tag_threadId,
  input  [3:0]  io_in_2_bits_tag_id,
  output        io_in_3_ready,
  input         io_in_3_valid,
  input  [63:0] io_in_3_bits_value,
  input         io_in_3_bits_isError,
  input         io_in_3_bits_tag_threadId,
  input  [3:0]  io_in_3_bits_tag_id,
  input         io_out_ready,
  output        io_out_valid,
  output        io_out_bits_resultType,
  output [63:0] io_out_bits_value,
  output        io_out_bits_isError,
  output        io_out_bits_tag_threadId,
  output [3:0]  io_out_bits_tag_id
);
  wire [63:0] _GEN_2 = io_in_2_valid ? io_in_2_bits_value : io_in_3_bits_value; // @[Arbiter.scala 136:15 138:26 140:19]
  wire  _GEN_3 = io_in_2_valid ? io_in_2_bits_isError : io_in_3_bits_isError; // @[Arbiter.scala 136:15 138:26 140:19]
  wire  _GEN_4 = io_in_2_valid ? io_in_2_bits_tag_threadId : io_in_3_bits_tag_threadId; // @[Arbiter.scala 136:15 138:26 140:19]
  wire [3:0] _GEN_5 = io_in_2_valid ? io_in_2_bits_tag_id : io_in_3_bits_tag_id; // @[Arbiter.scala 136:15 138:26 140:19]
  wire [63:0] _GEN_8 = io_in_1_valid ? io_in_1_bits_value : _GEN_2; // @[Arbiter.scala 138:26 140:19]
  wire  _GEN_9 = io_in_1_valid ? 1'h0 : _GEN_3; // @[Arbiter.scala 138:26 140:19]
  wire  _GEN_10 = io_in_1_valid ? io_in_1_bits_tag_threadId : _GEN_4; // @[Arbiter.scala 138:26 140:19]
  wire [3:0] _GEN_11 = io_in_1_valid ? io_in_1_bits_tag_id : _GEN_5; // @[Arbiter.scala 138:26 140:19]
  wire  grant_1 = ~io_in_0_valid; // @[Arbiter.scala 45:78]
  wire  grant_2 = ~(io_in_0_valid | io_in_1_valid); // @[Arbiter.scala 45:78]
  wire  grant_3 = ~(io_in_0_valid | io_in_1_valid | io_in_2_valid); // @[Arbiter.scala 45:78]
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 146:19]
  assign io_in_1_ready = grant_1 & io_out_ready; // @[Arbiter.scala 146:19]
  assign io_in_2_ready = grant_2 & io_out_ready; // @[Arbiter.scala 146:19]
  assign io_in_3_ready = grant_3 & io_out_ready; // @[Arbiter.scala 146:19]
  assign io_out_valid = ~grant_3 | io_in_3_valid; // @[Arbiter.scala 147:31]
  assign io_out_bits_resultType = io_in_0_valid ? io_in_0_bits_resultType : io_in_1_valid & io_in_1_bits_resultType; // @[Arbiter.scala 138:26 140:19]
  assign io_out_bits_value = io_in_0_valid ? io_in_0_bits_value : _GEN_8; // @[Arbiter.scala 138:26 140:19]
  assign io_out_bits_isError = io_in_0_valid ? 1'h0 : _GEN_9; // @[Arbiter.scala 138:26 140:19]
  assign io_out_bits_tag_threadId = io_in_0_valid ? io_in_0_bits_tag_threadId : _GEN_10; // @[Arbiter.scala 138:26 140:19]
  assign io_out_bits_tag_id = io_in_0_valid ? io_in_0_bits_tag_id : _GEN_11; // @[Arbiter.scala 138:26 140:19]
endmodule
module OutputCollector(
  input         clock,
  input         reset,
  output        io_outputs_0_outputs_valid,
  output        io_outputs_0_outputs_bits_resultType,
  output [63:0] io_outputs_0_outputs_bits_value,
  output        io_outputs_0_outputs_bits_isError,
  output        io_outputs_0_outputs_bits_tag_threadId,
  output [3:0]  io_outputs_0_outputs_bits_tag_id,
  output        io_outputs_1_outputs_valid,
  output        io_outputs_1_outputs_bits_resultType,
  output [63:0] io_outputs_1_outputs_bits_value,
  output        io_outputs_1_outputs_bits_isError,
  output        io_outputs_1_outputs_bits_tag_threadId,
  output [3:0]  io_outputs_1_outputs_bits_tag_id,
  output        io_executor_0_ready,
  input         io_executor_0_valid,
  input         io_executor_0_bits_resultType,
  input  [63:0] io_executor_0_bits_value,
  input         io_executor_0_bits_tag_threadId,
  input  [3:0]  io_executor_0_bits_tag_id,
  output        io_executor_1_ready,
  input         io_executor_1_valid,
  input         io_executor_1_bits_resultType,
  input  [63:0] io_executor_1_bits_value,
  input         io_executor_1_bits_tag_threadId,
  input  [3:0]  io_executor_1_bits_tag_id,
  output        io_dataMemory_ready,
  input         io_dataMemory_valid,
  input  [63:0] io_dataMemory_bits_value,
  input         io_dataMemory_bits_isError,
  input         io_dataMemory_bits_tag_threadId,
  input  [3:0]  io_dataMemory_bits_tag_id,
  output        io_csr_0_ready,
  input         io_csr_0_valid,
  input  [63:0] io_csr_0_bits_value,
  input         io_csr_0_bits_isError,
  input         io_csr_0_bits_tag_threadId,
  input  [3:0]  io_csr_0_bits_tag_id,
  output        io_csr_1_ready,
  input         io_csr_1_valid,
  input  [63:0] io_csr_1_bits_value,
  input         io_csr_1_bits_isError,
  input         io_csr_1_bits_tag_threadId,
  input  [3:0]  io_csr_1_bits_tag_id,
  input         io_isError_0,
  input         io_isError_1
);
  wire  threadsOutputQueue_0_clock; // @[OutputCollector.scala 20:36]
  wire  threadsOutputQueue_0_reset; // @[OutputCollector.scala 20:36]
  wire  threadsOutputQueue_0_input_ready; // @[OutputCollector.scala 20:36]
  wire  threadsOutputQueue_0_input_valid; // @[OutputCollector.scala 20:36]
  wire  threadsOutputQueue_0_input_bits_resultType; // @[OutputCollector.scala 20:36]
  wire [63:0] threadsOutputQueue_0_input_bits_value; // @[OutputCollector.scala 20:36]
  wire  threadsOutputQueue_0_input_bits_isError; // @[OutputCollector.scala 20:36]
  wire  threadsOutputQueue_0_input_bits_tag_threadId; // @[OutputCollector.scala 20:36]
  wire [3:0] threadsOutputQueue_0_input_bits_tag_id; // @[OutputCollector.scala 20:36]
  wire  threadsOutputQueue_0_output_valid; // @[OutputCollector.scala 20:36]
  wire  threadsOutputQueue_0_output_bits_resultType; // @[OutputCollector.scala 20:36]
  wire [63:0] threadsOutputQueue_0_output_bits_value; // @[OutputCollector.scala 20:36]
  wire  threadsOutputQueue_0_output_bits_isError; // @[OutputCollector.scala 20:36]
  wire  threadsOutputQueue_0_output_bits_tag_threadId; // @[OutputCollector.scala 20:36]
  wire [3:0] threadsOutputQueue_0_output_bits_tag_id; // @[OutputCollector.scala 20:36]
  wire  threadsOutputQueue_0_flush; // @[OutputCollector.scala 20:36]
  wire  threadsOutputQueue_1_clock; // @[OutputCollector.scala 20:36]
  wire  threadsOutputQueue_1_reset; // @[OutputCollector.scala 20:36]
  wire  threadsOutputQueue_1_input_ready; // @[OutputCollector.scala 20:36]
  wire  threadsOutputQueue_1_input_valid; // @[OutputCollector.scala 20:36]
  wire  threadsOutputQueue_1_input_bits_resultType; // @[OutputCollector.scala 20:36]
  wire [63:0] threadsOutputQueue_1_input_bits_value; // @[OutputCollector.scala 20:36]
  wire  threadsOutputQueue_1_input_bits_isError; // @[OutputCollector.scala 20:36]
  wire  threadsOutputQueue_1_input_bits_tag_threadId; // @[OutputCollector.scala 20:36]
  wire [3:0] threadsOutputQueue_1_input_bits_tag_id; // @[OutputCollector.scala 20:36]
  wire  threadsOutputQueue_1_output_valid; // @[OutputCollector.scala 20:36]
  wire  threadsOutputQueue_1_output_bits_resultType; // @[OutputCollector.scala 20:36]
  wire [63:0] threadsOutputQueue_1_output_bits_value; // @[OutputCollector.scala 20:36]
  wire  threadsOutputQueue_1_output_bits_isError; // @[OutputCollector.scala 20:36]
  wire  threadsOutputQueue_1_output_bits_tag_threadId; // @[OutputCollector.scala 20:36]
  wire [3:0] threadsOutputQueue_1_output_bits_tag_id; // @[OutputCollector.scala 20:36]
  wire  threadsOutputQueue_1_flush; // @[OutputCollector.scala 20:36]
  wire  threadsArbiter_0_io_in_0_ready; // @[OutputCollector.scala 23:13]
  wire  threadsArbiter_0_io_in_0_valid; // @[OutputCollector.scala 23:13]
  wire  threadsArbiter_0_io_in_0_bits_resultType; // @[OutputCollector.scala 23:13]
  wire [63:0] threadsArbiter_0_io_in_0_bits_value; // @[OutputCollector.scala 23:13]
  wire  threadsArbiter_0_io_in_0_bits_tag_threadId; // @[OutputCollector.scala 23:13]
  wire [3:0] threadsArbiter_0_io_in_0_bits_tag_id; // @[OutputCollector.scala 23:13]
  wire  threadsArbiter_0_io_in_1_ready; // @[OutputCollector.scala 23:13]
  wire  threadsArbiter_0_io_in_1_valid; // @[OutputCollector.scala 23:13]
  wire  threadsArbiter_0_io_in_1_bits_resultType; // @[OutputCollector.scala 23:13]
  wire [63:0] threadsArbiter_0_io_in_1_bits_value; // @[OutputCollector.scala 23:13]
  wire  threadsArbiter_0_io_in_1_bits_tag_threadId; // @[OutputCollector.scala 23:13]
  wire [3:0] threadsArbiter_0_io_in_1_bits_tag_id; // @[OutputCollector.scala 23:13]
  wire  threadsArbiter_0_io_in_2_ready; // @[OutputCollector.scala 23:13]
  wire  threadsArbiter_0_io_in_2_valid; // @[OutputCollector.scala 23:13]
  wire [63:0] threadsArbiter_0_io_in_2_bits_value; // @[OutputCollector.scala 23:13]
  wire  threadsArbiter_0_io_in_2_bits_isError; // @[OutputCollector.scala 23:13]
  wire  threadsArbiter_0_io_in_2_bits_tag_threadId; // @[OutputCollector.scala 23:13]
  wire [3:0] threadsArbiter_0_io_in_2_bits_tag_id; // @[OutputCollector.scala 23:13]
  wire  threadsArbiter_0_io_in_3_ready; // @[OutputCollector.scala 23:13]
  wire  threadsArbiter_0_io_in_3_valid; // @[OutputCollector.scala 23:13]
  wire [63:0] threadsArbiter_0_io_in_3_bits_value; // @[OutputCollector.scala 23:13]
  wire  threadsArbiter_0_io_in_3_bits_isError; // @[OutputCollector.scala 23:13]
  wire  threadsArbiter_0_io_in_3_bits_tag_threadId; // @[OutputCollector.scala 23:13]
  wire [3:0] threadsArbiter_0_io_in_3_bits_tag_id; // @[OutputCollector.scala 23:13]
  wire  threadsArbiter_0_io_out_ready; // @[OutputCollector.scala 23:13]
  wire  threadsArbiter_0_io_out_valid; // @[OutputCollector.scala 23:13]
  wire  threadsArbiter_0_io_out_bits_resultType; // @[OutputCollector.scala 23:13]
  wire [63:0] threadsArbiter_0_io_out_bits_value; // @[OutputCollector.scala 23:13]
  wire  threadsArbiter_0_io_out_bits_isError; // @[OutputCollector.scala 23:13]
  wire  threadsArbiter_0_io_out_bits_tag_threadId; // @[OutputCollector.scala 23:13]
  wire [3:0] threadsArbiter_0_io_out_bits_tag_id; // @[OutputCollector.scala 23:13]
  wire  threadsArbiter_1_io_in_0_ready; // @[OutputCollector.scala 23:13]
  wire  threadsArbiter_1_io_in_0_valid; // @[OutputCollector.scala 23:13]
  wire  threadsArbiter_1_io_in_0_bits_resultType; // @[OutputCollector.scala 23:13]
  wire [63:0] threadsArbiter_1_io_in_0_bits_value; // @[OutputCollector.scala 23:13]
  wire  threadsArbiter_1_io_in_0_bits_tag_threadId; // @[OutputCollector.scala 23:13]
  wire [3:0] threadsArbiter_1_io_in_0_bits_tag_id; // @[OutputCollector.scala 23:13]
  wire  threadsArbiter_1_io_in_1_ready; // @[OutputCollector.scala 23:13]
  wire  threadsArbiter_1_io_in_1_valid; // @[OutputCollector.scala 23:13]
  wire  threadsArbiter_1_io_in_1_bits_resultType; // @[OutputCollector.scala 23:13]
  wire [63:0] threadsArbiter_1_io_in_1_bits_value; // @[OutputCollector.scala 23:13]
  wire  threadsArbiter_1_io_in_1_bits_tag_threadId; // @[OutputCollector.scala 23:13]
  wire [3:0] threadsArbiter_1_io_in_1_bits_tag_id; // @[OutputCollector.scala 23:13]
  wire  threadsArbiter_1_io_in_2_ready; // @[OutputCollector.scala 23:13]
  wire  threadsArbiter_1_io_in_2_valid; // @[OutputCollector.scala 23:13]
  wire [63:0] threadsArbiter_1_io_in_2_bits_value; // @[OutputCollector.scala 23:13]
  wire  threadsArbiter_1_io_in_2_bits_isError; // @[OutputCollector.scala 23:13]
  wire  threadsArbiter_1_io_in_2_bits_tag_threadId; // @[OutputCollector.scala 23:13]
  wire [3:0] threadsArbiter_1_io_in_2_bits_tag_id; // @[OutputCollector.scala 23:13]
  wire  threadsArbiter_1_io_in_3_ready; // @[OutputCollector.scala 23:13]
  wire  threadsArbiter_1_io_in_3_valid; // @[OutputCollector.scala 23:13]
  wire [63:0] threadsArbiter_1_io_in_3_bits_value; // @[OutputCollector.scala 23:13]
  wire  threadsArbiter_1_io_in_3_bits_isError; // @[OutputCollector.scala 23:13]
  wire  threadsArbiter_1_io_in_3_bits_tag_threadId; // @[OutputCollector.scala 23:13]
  wire [3:0] threadsArbiter_1_io_in_3_bits_tag_id; // @[OutputCollector.scala 23:13]
  wire  threadsArbiter_1_io_out_ready; // @[OutputCollector.scala 23:13]
  wire  threadsArbiter_1_io_out_valid; // @[OutputCollector.scala 23:13]
  wire  threadsArbiter_1_io_out_bits_resultType; // @[OutputCollector.scala 23:13]
  wire [63:0] threadsArbiter_1_io_out_bits_value; // @[OutputCollector.scala 23:13]
  wire  threadsArbiter_1_io_out_bits_isError; // @[OutputCollector.scala 23:13]
  wire  threadsArbiter_1_io_out_bits_tag_threadId; // @[OutputCollector.scala 23:13]
  wire [3:0] threadsArbiter_1_io_out_bits_tag_id; // @[OutputCollector.scala 23:13]
  wire  _threadsArbiter_0_io_in_0_valid_T = ~io_executor_0_bits_tag_threadId; // @[OutputCollector.scala 33:52]
  wire  _threadsArbiter_0_io_in_1_valid_T = ~io_executor_1_bits_tag_threadId; // @[OutputCollector.scala 33:52]
  wire  _threadsArbiter_0_io_in_2_valid_T = ~io_dataMemory_bits_tag_threadId; // @[OutputCollector.scala 38:72]
  wire  _io_executor_0_ready_T_1 = threadsArbiter_0_io_in_0_ready & _threadsArbiter_0_io_in_0_valid_T; // @[OutputCollector.scala 50:18]
  wire  _io_executor_0_ready_T_3 = threadsArbiter_1_io_in_0_ready & io_executor_0_bits_tag_threadId; // @[OutputCollector.scala 50:18]
  wire  _io_executor_1_ready_T_1 = threadsArbiter_0_io_in_1_ready & _threadsArbiter_0_io_in_1_valid_T; // @[OutputCollector.scala 50:18]
  wire  _io_executor_1_ready_T_3 = threadsArbiter_1_io_in_1_ready & io_executor_1_bits_tag_threadId; // @[OutputCollector.scala 50:18]
  wire  _io_dataMemory_ready_T_1 = threadsArbiter_0_io_in_2_ready & _threadsArbiter_0_io_in_2_valid_T; // @[OutputCollector.scala 58:16]
  wire  _io_dataMemory_ready_T_3 = threadsArbiter_1_io_in_2_ready & io_dataMemory_bits_tag_threadId; // @[OutputCollector.scala 58:16]
  FIFO_1 threadsOutputQueue_0 ( // @[OutputCollector.scala 20:36]
    .clock(threadsOutputQueue_0_clock),
    .reset(threadsOutputQueue_0_reset),
    .input_ready(threadsOutputQueue_0_input_ready),
    .input_valid(threadsOutputQueue_0_input_valid),
    .input_bits_resultType(threadsOutputQueue_0_input_bits_resultType),
    .input_bits_value(threadsOutputQueue_0_input_bits_value),
    .input_bits_isError(threadsOutputQueue_0_input_bits_isError),
    .input_bits_tag_threadId(threadsOutputQueue_0_input_bits_tag_threadId),
    .input_bits_tag_id(threadsOutputQueue_0_input_bits_tag_id),
    .output_valid(threadsOutputQueue_0_output_valid),
    .output_bits_resultType(threadsOutputQueue_0_output_bits_resultType),
    .output_bits_value(threadsOutputQueue_0_output_bits_value),
    .output_bits_isError(threadsOutputQueue_0_output_bits_isError),
    .output_bits_tag_threadId(threadsOutputQueue_0_output_bits_tag_threadId),
    .output_bits_tag_id(threadsOutputQueue_0_output_bits_tag_id),
    .flush(threadsOutputQueue_0_flush)
  );
  FIFO_1 threadsOutputQueue_1 ( // @[OutputCollector.scala 20:36]
    .clock(threadsOutputQueue_1_clock),
    .reset(threadsOutputQueue_1_reset),
    .input_ready(threadsOutputQueue_1_input_ready),
    .input_valid(threadsOutputQueue_1_input_valid),
    .input_bits_resultType(threadsOutputQueue_1_input_bits_resultType),
    .input_bits_value(threadsOutputQueue_1_input_bits_value),
    .input_bits_isError(threadsOutputQueue_1_input_bits_isError),
    .input_bits_tag_threadId(threadsOutputQueue_1_input_bits_tag_threadId),
    .input_bits_tag_id(threadsOutputQueue_1_input_bits_tag_id),
    .output_valid(threadsOutputQueue_1_output_valid),
    .output_bits_resultType(threadsOutputQueue_1_output_bits_resultType),
    .output_bits_value(threadsOutputQueue_1_output_bits_value),
    .output_bits_isError(threadsOutputQueue_1_output_bits_isError),
    .output_bits_tag_threadId(threadsOutputQueue_1_output_bits_tag_threadId),
    .output_bits_tag_id(threadsOutputQueue_1_output_bits_tag_id),
    .flush(threadsOutputQueue_1_flush)
  );
  Arbiter threadsArbiter_0 ( // @[OutputCollector.scala 23:13]
    .io_in_0_ready(threadsArbiter_0_io_in_0_ready),
    .io_in_0_valid(threadsArbiter_0_io_in_0_valid),
    .io_in_0_bits_resultType(threadsArbiter_0_io_in_0_bits_resultType),
    .io_in_0_bits_value(threadsArbiter_0_io_in_0_bits_value),
    .io_in_0_bits_tag_threadId(threadsArbiter_0_io_in_0_bits_tag_threadId),
    .io_in_0_bits_tag_id(threadsArbiter_0_io_in_0_bits_tag_id),
    .io_in_1_ready(threadsArbiter_0_io_in_1_ready),
    .io_in_1_valid(threadsArbiter_0_io_in_1_valid),
    .io_in_1_bits_resultType(threadsArbiter_0_io_in_1_bits_resultType),
    .io_in_1_bits_value(threadsArbiter_0_io_in_1_bits_value),
    .io_in_1_bits_tag_threadId(threadsArbiter_0_io_in_1_bits_tag_threadId),
    .io_in_1_bits_tag_id(threadsArbiter_0_io_in_1_bits_tag_id),
    .io_in_2_ready(threadsArbiter_0_io_in_2_ready),
    .io_in_2_valid(threadsArbiter_0_io_in_2_valid),
    .io_in_2_bits_value(threadsArbiter_0_io_in_2_bits_value),
    .io_in_2_bits_isError(threadsArbiter_0_io_in_2_bits_isError),
    .io_in_2_bits_tag_threadId(threadsArbiter_0_io_in_2_bits_tag_threadId),
    .io_in_2_bits_tag_id(threadsArbiter_0_io_in_2_bits_tag_id),
    .io_in_3_ready(threadsArbiter_0_io_in_3_ready),
    .io_in_3_valid(threadsArbiter_0_io_in_3_valid),
    .io_in_3_bits_value(threadsArbiter_0_io_in_3_bits_value),
    .io_in_3_bits_isError(threadsArbiter_0_io_in_3_bits_isError),
    .io_in_3_bits_tag_threadId(threadsArbiter_0_io_in_3_bits_tag_threadId),
    .io_in_3_bits_tag_id(threadsArbiter_0_io_in_3_bits_tag_id),
    .io_out_ready(threadsArbiter_0_io_out_ready),
    .io_out_valid(threadsArbiter_0_io_out_valid),
    .io_out_bits_resultType(threadsArbiter_0_io_out_bits_resultType),
    .io_out_bits_value(threadsArbiter_0_io_out_bits_value),
    .io_out_bits_isError(threadsArbiter_0_io_out_bits_isError),
    .io_out_bits_tag_threadId(threadsArbiter_0_io_out_bits_tag_threadId),
    .io_out_bits_tag_id(threadsArbiter_0_io_out_bits_tag_id)
  );
  Arbiter threadsArbiter_1 ( // @[OutputCollector.scala 23:13]
    .io_in_0_ready(threadsArbiter_1_io_in_0_ready),
    .io_in_0_valid(threadsArbiter_1_io_in_0_valid),
    .io_in_0_bits_resultType(threadsArbiter_1_io_in_0_bits_resultType),
    .io_in_0_bits_value(threadsArbiter_1_io_in_0_bits_value),
    .io_in_0_bits_tag_threadId(threadsArbiter_1_io_in_0_bits_tag_threadId),
    .io_in_0_bits_tag_id(threadsArbiter_1_io_in_0_bits_tag_id),
    .io_in_1_ready(threadsArbiter_1_io_in_1_ready),
    .io_in_1_valid(threadsArbiter_1_io_in_1_valid),
    .io_in_1_bits_resultType(threadsArbiter_1_io_in_1_bits_resultType),
    .io_in_1_bits_value(threadsArbiter_1_io_in_1_bits_value),
    .io_in_1_bits_tag_threadId(threadsArbiter_1_io_in_1_bits_tag_threadId),
    .io_in_1_bits_tag_id(threadsArbiter_1_io_in_1_bits_tag_id),
    .io_in_2_ready(threadsArbiter_1_io_in_2_ready),
    .io_in_2_valid(threadsArbiter_1_io_in_2_valid),
    .io_in_2_bits_value(threadsArbiter_1_io_in_2_bits_value),
    .io_in_2_bits_isError(threadsArbiter_1_io_in_2_bits_isError),
    .io_in_2_bits_tag_threadId(threadsArbiter_1_io_in_2_bits_tag_threadId),
    .io_in_2_bits_tag_id(threadsArbiter_1_io_in_2_bits_tag_id),
    .io_in_3_ready(threadsArbiter_1_io_in_3_ready),
    .io_in_3_valid(threadsArbiter_1_io_in_3_valid),
    .io_in_3_bits_value(threadsArbiter_1_io_in_3_bits_value),
    .io_in_3_bits_isError(threadsArbiter_1_io_in_3_bits_isError),
    .io_in_3_bits_tag_threadId(threadsArbiter_1_io_in_3_bits_tag_threadId),
    .io_in_3_bits_tag_id(threadsArbiter_1_io_in_3_bits_tag_id),
    .io_out_ready(threadsArbiter_1_io_out_ready),
    .io_out_valid(threadsArbiter_1_io_out_valid),
    .io_out_bits_resultType(threadsArbiter_1_io_out_bits_resultType),
    .io_out_bits_value(threadsArbiter_1_io_out_bits_value),
    .io_out_bits_isError(threadsArbiter_1_io_out_bits_isError),
    .io_out_bits_tag_threadId(threadsArbiter_1_io_out_bits_tag_threadId),
    .io_out_bits_tag_id(threadsArbiter_1_io_out_bits_tag_id)
  );
  assign io_outputs_0_outputs_valid = threadsOutputQueue_0_output_valid; // @[OutputCollector.scala 63:33]
  assign io_outputs_0_outputs_bits_resultType = threadsOutputQueue_0_output_bits_resultType; // @[OutputCollector.scala 64:32]
  assign io_outputs_0_outputs_bits_value = threadsOutputQueue_0_output_bits_value; // @[OutputCollector.scala 64:32]
  assign io_outputs_0_outputs_bits_isError = threadsOutputQueue_0_output_bits_isError; // @[OutputCollector.scala 64:32]
  assign io_outputs_0_outputs_bits_tag_threadId = threadsOutputQueue_0_output_bits_tag_threadId; // @[OutputCollector.scala 64:32]
  assign io_outputs_0_outputs_bits_tag_id = threadsOutputQueue_0_output_bits_tag_id; // @[OutputCollector.scala 64:32]
  assign io_outputs_1_outputs_valid = threadsOutputQueue_1_output_valid; // @[OutputCollector.scala 63:33]
  assign io_outputs_1_outputs_bits_resultType = threadsOutputQueue_1_output_bits_resultType; // @[OutputCollector.scala 64:32]
  assign io_outputs_1_outputs_bits_value = threadsOutputQueue_1_output_bits_value; // @[OutputCollector.scala 64:32]
  assign io_outputs_1_outputs_bits_isError = threadsOutputQueue_1_output_bits_isError; // @[OutputCollector.scala 64:32]
  assign io_outputs_1_outputs_bits_tag_threadId = threadsOutputQueue_1_output_bits_tag_threadId; // @[OutputCollector.scala 64:32]
  assign io_outputs_1_outputs_bits_tag_id = threadsOutputQueue_1_output_bits_tag_id; // @[OutputCollector.scala 64:32]
  assign io_executor_0_ready = _io_executor_0_ready_T_1 | _io_executor_0_ready_T_3; // @[OutputCollector.scala 52:17]
  assign io_executor_1_ready = _io_executor_1_ready_T_1 | _io_executor_1_ready_T_3; // @[OutputCollector.scala 52:17]
  assign io_dataMemory_ready = _io_dataMemory_ready_T_1 | _io_dataMemory_ready_T_3; // @[OutputCollector.scala 60:15]
  assign io_csr_0_ready = threadsArbiter_0_io_in_3_ready; // @[OutputCollector.scala 39:53]
  assign io_csr_1_ready = threadsArbiter_1_io_in_3_ready; // @[OutputCollector.scala 39:53]
  assign threadsOutputQueue_0_clock = clock;
  assign threadsOutputQueue_0_reset = reset;
  assign threadsOutputQueue_0_input_valid = threadsArbiter_0_io_out_valid; // @[OutputCollector.scala 41:35]
  assign threadsOutputQueue_0_input_bits_resultType = threadsArbiter_0_io_out_bits_resultType; // @[OutputCollector.scala 41:35]
  assign threadsOutputQueue_0_input_bits_value = threadsArbiter_0_io_out_bits_value; // @[OutputCollector.scala 41:35]
  assign threadsOutputQueue_0_input_bits_isError = threadsArbiter_0_io_out_bits_isError; // @[OutputCollector.scala 41:35]
  assign threadsOutputQueue_0_input_bits_tag_threadId = threadsArbiter_0_io_out_bits_tag_threadId; // @[OutputCollector.scala 41:35]
  assign threadsOutputQueue_0_input_bits_tag_id = threadsArbiter_0_io_out_bits_tag_id; // @[OutputCollector.scala 41:35]
  assign threadsOutputQueue_0_flush = io_isError_0; // @[OutputCollector.scala 42:35]
  assign threadsOutputQueue_1_clock = clock;
  assign threadsOutputQueue_1_reset = reset;
  assign threadsOutputQueue_1_input_valid = threadsArbiter_1_io_out_valid; // @[OutputCollector.scala 41:35]
  assign threadsOutputQueue_1_input_bits_resultType = threadsArbiter_1_io_out_bits_resultType; // @[OutputCollector.scala 41:35]
  assign threadsOutputQueue_1_input_bits_value = threadsArbiter_1_io_out_bits_value; // @[OutputCollector.scala 41:35]
  assign threadsOutputQueue_1_input_bits_isError = threadsArbiter_1_io_out_bits_isError; // @[OutputCollector.scala 41:35]
  assign threadsOutputQueue_1_input_bits_tag_threadId = threadsArbiter_1_io_out_bits_tag_threadId; // @[OutputCollector.scala 41:35]
  assign threadsOutputQueue_1_input_bits_tag_id = threadsArbiter_1_io_out_bits_tag_id; // @[OutputCollector.scala 41:35]
  assign threadsOutputQueue_1_flush = io_isError_1; // @[OutputCollector.scala 42:35]
  assign threadsArbiter_0_io_in_0_valid = io_executor_0_valid & ~io_executor_0_bits_tag_threadId; // @[OutputCollector.scala 33:16]
  assign threadsArbiter_0_io_in_0_bits_resultType = io_executor_0_bits_resultType; // @[OutputCollector.scala 28:36]
  assign threadsArbiter_0_io_in_0_bits_value = io_executor_0_bits_value; // @[OutputCollector.scala 28:36]
  assign threadsArbiter_0_io_in_0_bits_tag_threadId = io_executor_0_bits_tag_threadId; // @[OutputCollector.scala 28:36]
  assign threadsArbiter_0_io_in_0_bits_tag_id = io_executor_0_bits_tag_id; // @[OutputCollector.scala 28:36]
  assign threadsArbiter_0_io_in_1_valid = io_executor_1_valid & ~io_executor_1_bits_tag_threadId; // @[OutputCollector.scala 33:16]
  assign threadsArbiter_0_io_in_1_bits_resultType = io_executor_1_bits_resultType; // @[OutputCollector.scala 28:36]
  assign threadsArbiter_0_io_in_1_bits_value = io_executor_1_bits_value; // @[OutputCollector.scala 28:36]
  assign threadsArbiter_0_io_in_1_bits_tag_threadId = io_executor_1_bits_tag_threadId; // @[OutputCollector.scala 28:36]
  assign threadsArbiter_0_io_in_1_bits_tag_id = io_executor_1_bits_tag_id; // @[OutputCollector.scala 28:36]
  assign threadsArbiter_0_io_in_2_valid = io_dataMemory_valid & ~io_dataMemory_bits_tag_threadId; // @[OutputCollector.scala 38:37]
  assign threadsArbiter_0_io_in_2_bits_value = io_dataMemory_bits_value; // @[OutputCollector.scala 35:49]
  assign threadsArbiter_0_io_in_2_bits_isError = io_dataMemory_bits_isError; // @[OutputCollector.scala 35:49]
  assign threadsArbiter_0_io_in_2_bits_tag_threadId = io_dataMemory_bits_tag_threadId; // @[OutputCollector.scala 35:49]
  assign threadsArbiter_0_io_in_2_bits_tag_id = io_dataMemory_bits_tag_id; // @[OutputCollector.scala 35:49]
  assign threadsArbiter_0_io_in_3_valid = io_csr_0_valid; // @[OutputCollector.scala 39:53]
  assign threadsArbiter_0_io_in_3_bits_value = io_csr_0_bits_value; // @[OutputCollector.scala 39:53]
  assign threadsArbiter_0_io_in_3_bits_isError = io_csr_0_bits_isError; // @[OutputCollector.scala 39:53]
  assign threadsArbiter_0_io_in_3_bits_tag_threadId = io_csr_0_bits_tag_threadId; // @[OutputCollector.scala 39:53]
  assign threadsArbiter_0_io_in_3_bits_tag_id = io_csr_0_bits_tag_id; // @[OutputCollector.scala 39:53]
  assign threadsArbiter_0_io_out_ready = threadsOutputQueue_0_input_ready; // @[OutputCollector.scala 41:35]
  assign threadsArbiter_1_io_in_0_valid = io_executor_0_valid & io_executor_0_bits_tag_threadId; // @[OutputCollector.scala 33:16]
  assign threadsArbiter_1_io_in_0_bits_resultType = io_executor_0_bits_resultType; // @[OutputCollector.scala 28:36]
  assign threadsArbiter_1_io_in_0_bits_value = io_executor_0_bits_value; // @[OutputCollector.scala 28:36]
  assign threadsArbiter_1_io_in_0_bits_tag_threadId = io_executor_0_bits_tag_threadId; // @[OutputCollector.scala 28:36]
  assign threadsArbiter_1_io_in_0_bits_tag_id = io_executor_0_bits_tag_id; // @[OutputCollector.scala 28:36]
  assign threadsArbiter_1_io_in_1_valid = io_executor_1_valid & io_executor_1_bits_tag_threadId; // @[OutputCollector.scala 33:16]
  assign threadsArbiter_1_io_in_1_bits_resultType = io_executor_1_bits_resultType; // @[OutputCollector.scala 28:36]
  assign threadsArbiter_1_io_in_1_bits_value = io_executor_1_bits_value; // @[OutputCollector.scala 28:36]
  assign threadsArbiter_1_io_in_1_bits_tag_threadId = io_executor_1_bits_tag_threadId; // @[OutputCollector.scala 28:36]
  assign threadsArbiter_1_io_in_1_bits_tag_id = io_executor_1_bits_tag_id; // @[OutputCollector.scala 28:36]
  assign threadsArbiter_1_io_in_2_valid = io_dataMemory_valid & io_dataMemory_bits_tag_threadId; // @[OutputCollector.scala 38:37]
  assign threadsArbiter_1_io_in_2_bits_value = io_dataMemory_bits_value; // @[OutputCollector.scala 35:49]
  assign threadsArbiter_1_io_in_2_bits_isError = io_dataMemory_bits_isError; // @[OutputCollector.scala 35:49]
  assign threadsArbiter_1_io_in_2_bits_tag_threadId = io_dataMemory_bits_tag_threadId; // @[OutputCollector.scala 35:49]
  assign threadsArbiter_1_io_in_2_bits_tag_id = io_dataMemory_bits_tag_id; // @[OutputCollector.scala 35:49]
  assign threadsArbiter_1_io_in_3_valid = io_csr_1_valid; // @[OutputCollector.scala 39:53]
  assign threadsArbiter_1_io_in_3_bits_value = io_csr_1_bits_value; // @[OutputCollector.scala 39:53]
  assign threadsArbiter_1_io_in_3_bits_isError = io_csr_1_bits_isError; // @[OutputCollector.scala 39:53]
  assign threadsArbiter_1_io_in_3_bits_tag_threadId = io_csr_1_bits_tag_threadId; // @[OutputCollector.scala 39:53]
  assign threadsArbiter_1_io_in_3_bits_tag_id = io_csr_1_bits_tag_id; // @[OutputCollector.scala 39:53]
  assign threadsArbiter_1_io_out_ready = threadsOutputQueue_1_input_ready; // @[OutputCollector.scala 41:35]
endmodule
module Queue_3(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input         io_enq_bits_threadId,
  input  [63:0] io_enq_bits_programCounterOffset,
  output        io_deq_valid,
  output        io_deq_bits_threadId,
  output [63:0] io_deq_bits_programCounterOffset,
  input         io_flush
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_3;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  reg  ram_threadId [0:3]; // @[Decoupled.scala 273:44]
  wire  ram_threadId_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:44]
  wire [1:0] ram_threadId_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:44]
  wire  ram_threadId_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:44]
  wire  ram_threadId_MPORT_data; // @[Decoupled.scala 273:44]
  wire [1:0] ram_threadId_MPORT_addr; // @[Decoupled.scala 273:44]
  wire  ram_threadId_MPORT_mask; // @[Decoupled.scala 273:44]
  wire  ram_threadId_MPORT_en; // @[Decoupled.scala 273:44]
  reg  ram_threadId_io_deq_bits_MPORT_en_pipe_0;
  reg [1:0] ram_threadId_io_deq_bits_MPORT_addr_pipe_0;
  reg [63:0] ram_programCounterOffset [0:3]; // @[Decoupled.scala 273:44]
  wire  ram_programCounterOffset_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:44]
  wire [1:0] ram_programCounterOffset_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:44]
  wire [63:0] ram_programCounterOffset_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:44]
  wire [63:0] ram_programCounterOffset_MPORT_data; // @[Decoupled.scala 273:44]
  wire [1:0] ram_programCounterOffset_MPORT_addr; // @[Decoupled.scala 273:44]
  wire  ram_programCounterOffset_MPORT_mask; // @[Decoupled.scala 273:44]
  wire  ram_programCounterOffset_MPORT_en; // @[Decoupled.scala 273:44]
  reg  ram_programCounterOffset_io_deq_bits_MPORT_en_pipe_0;
  reg [1:0] ram_programCounterOffset_io_deq_bits_MPORT_addr_pipe_0;
  reg [1:0] enq_ptr_value; // @[Counter.scala 61:40]
  reg [1:0] deq_ptr_value; // @[Counter.scala 61:40]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 277:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 278:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 279:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire [1:0] _value_T_1 = enq_ptr_value + 2'h1; // @[Counter.scala 77:24]
  wire [1:0] _value_T_3 = deq_ptr_value + 2'h1; // @[Counter.scala 77:24]
  wire [2:0] _deq_ptr_next_T_1 = 3'h4 - 3'h1; // @[Decoupled.scala 306:57]
  wire [2:0] _GEN_16 = {{1'd0}, deq_ptr_value}; // @[Decoupled.scala 306:42]
  assign ram_threadId_io_deq_bits_MPORT_en = ram_threadId_io_deq_bits_MPORT_en_pipe_0;
  assign ram_threadId_io_deq_bits_MPORT_addr = ram_threadId_io_deq_bits_MPORT_addr_pipe_0;
  assign ram_threadId_io_deq_bits_MPORT_data = ram_threadId[ram_threadId_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:44]
  assign ram_threadId_MPORT_data = io_enq_bits_threadId;
  assign ram_threadId_MPORT_addr = enq_ptr_value;
  assign ram_threadId_MPORT_mask = 1'h1;
  assign ram_threadId_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_programCounterOffset_io_deq_bits_MPORT_en = ram_programCounterOffset_io_deq_bits_MPORT_en_pipe_0;
  assign ram_programCounterOffset_io_deq_bits_MPORT_addr = ram_programCounterOffset_io_deq_bits_MPORT_addr_pipe_0;
  assign ram_programCounterOffset_io_deq_bits_MPORT_data =
    ram_programCounterOffset[ram_programCounterOffset_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:44]
  assign ram_programCounterOffset_MPORT_data = io_enq_bits_programCounterOffset;
  assign ram_programCounterOffset_MPORT_addr = enq_ptr_value;
  assign ram_programCounterOffset_MPORT_mask = 1'h1;
  assign ram_programCounterOffset_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 303:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 302:19]
  assign io_deq_bits_threadId = ram_threadId_io_deq_bits_MPORT_data; // @[Decoupled.scala 308:17]
  assign io_deq_bits_programCounterOffset = ram_programCounterOffset_io_deq_bits_MPORT_data; // @[Decoupled.scala 308:17]
  always @(posedge clock) begin
    if (ram_threadId_MPORT_en & ram_threadId_MPORT_mask) begin
      ram_threadId[ram_threadId_MPORT_addr] <= ram_threadId_MPORT_data; // @[Decoupled.scala 273:44]
    end
    ram_threadId_io_deq_bits_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (io_deq_valid) begin
        if (_GEN_16 == _deq_ptr_next_T_1) begin // @[Decoupled.scala 306:27]
          ram_threadId_io_deq_bits_MPORT_addr_pipe_0 <= 2'h0;
        end else begin
          ram_threadId_io_deq_bits_MPORT_addr_pipe_0 <= _value_T_3;
        end
      end else begin
        ram_threadId_io_deq_bits_MPORT_addr_pipe_0 <= deq_ptr_value;
      end
    end
    if (ram_programCounterOffset_MPORT_en & ram_programCounterOffset_MPORT_mask) begin
      ram_programCounterOffset[ram_programCounterOffset_MPORT_addr] <= ram_programCounterOffset_MPORT_data; // @[Decoupled.scala 273:44]
    end
    ram_programCounterOffset_io_deq_bits_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (io_deq_valid) begin
        if (_GEN_16 == _deq_ptr_next_T_1) begin // @[Decoupled.scala 306:27]
          ram_programCounterOffset_io_deq_bits_MPORT_addr_pipe_0 <= 2'h0;
        end else begin
          ram_programCounterOffset_io_deq_bits_MPORT_addr_pipe_0 <= _value_T_3;
        end
      end else begin
        ram_programCounterOffset_io_deq_bits_MPORT_addr_pipe_0 <= deq_ptr_value;
      end
    end
    if (reset) begin // @[Counter.scala 61:40]
      enq_ptr_value <= 2'h0; // @[Counter.scala 61:40]
    end else if (io_flush) begin // @[Decoupled.scala 296:15]
      enq_ptr_value <= 2'h0; // @[Counter.scala 98:11]
    end else if (do_enq) begin // @[Decoupled.scala 286:16]
      enq_ptr_value <= _value_T_1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      deq_ptr_value <= 2'h0; // @[Counter.scala 61:40]
    end else if (io_flush) begin // @[Decoupled.scala 296:15]
      deq_ptr_value <= 2'h0; // @[Counter.scala 98:11]
    end else if (io_deq_valid) begin // @[Decoupled.scala 290:16]
      deq_ptr_value <= _value_T_3; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (io_flush) begin // @[Decoupled.scala 296:15]
      maybe_full <= 1'h0; // @[Decoupled.scala 299:16]
    end else if (do_enq != io_deq_valid) begin // @[Decoupled.scala 293:27]
      maybe_full <= do_enq; // @[Decoupled.scala 294:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_threadId[initvar] = _RAND_0[0:0];
  _RAND_3 = {2{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_programCounterOffset[initvar] = _RAND_3[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_threadId_io_deq_bits_MPORT_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  ram_threadId_io_deq_bits_MPORT_addr_pipe_0 = _RAND_2[1:0];
  _RAND_4 = {1{`RANDOM}};
  ram_programCounterOffset_io_deq_bits_MPORT_en_pipe_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  ram_programCounterOffset_io_deq_bits_MPORT_addr_pipe_0 = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  enq_ptr_value = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  deq_ptr_value = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  maybe_full = _RAND_8[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module FIFO_3(
  input         clock,
  input         reset,
  output        input_ready,
  input         input_valid,
  input         input_bits_threadId,
  input  [63:0] input_bits_programCounterOffset,
  output        output_valid,
  output        output_bits_threadId,
  output [63:0] output_bits_programCounterOffset,
  input         flush
);
  wire  queue_clock; // @[FIFO.scala 16:29]
  wire  queue_reset; // @[FIFO.scala 16:29]
  wire  queue_io_enq_ready; // @[FIFO.scala 16:29]
  wire  queue_io_enq_valid; // @[FIFO.scala 16:29]
  wire  queue_io_enq_bits_threadId; // @[FIFO.scala 16:29]
  wire [63:0] queue_io_enq_bits_programCounterOffset; // @[FIFO.scala 16:29]
  wire  queue_io_deq_valid; // @[FIFO.scala 16:29]
  wire  queue_io_deq_bits_threadId; // @[FIFO.scala 16:29]
  wire [63:0] queue_io_deq_bits_programCounterOffset; // @[FIFO.scala 16:29]
  wire  queue_io_flush; // @[FIFO.scala 16:29]
  Queue_3 queue ( // @[FIFO.scala 16:29]
    .clock(queue_clock),
    .reset(queue_reset),
    .io_enq_ready(queue_io_enq_ready),
    .io_enq_valid(queue_io_enq_valid),
    .io_enq_bits_threadId(queue_io_enq_bits_threadId),
    .io_enq_bits_programCounterOffset(queue_io_enq_bits_programCounterOffset),
    .io_deq_valid(queue_io_deq_valid),
    .io_deq_bits_threadId(queue_io_deq_bits_threadId),
    .io_deq_bits_programCounterOffset(queue_io_deq_bits_programCounterOffset),
    .io_flush(queue_io_flush)
  );
  assign input_ready = queue_io_enq_ready; // @[FIFO.scala 19:16]
  assign output_valid = queue_io_deq_valid; // @[FIFO.scala 20:10]
  assign output_bits_threadId = queue_io_deq_bits_threadId; // @[FIFO.scala 20:10]
  assign output_bits_programCounterOffset = queue_io_deq_bits_programCounterOffset; // @[FIFO.scala 20:10]
  assign queue_clock = clock;
  assign queue_reset = reset;
  assign queue_io_enq_valid = input_valid; // @[FIFO.scala 19:16]
  assign queue_io_enq_bits_threadId = input_bits_threadId; // @[FIFO.scala 19:16]
  assign queue_io_enq_bits_programCounterOffset = input_bits_programCounterOffset; // @[FIFO.scala 19:16]
  assign queue_io_flush = flush; // @[FIFO.scala 23:15]
endmodule
module Arbiter_2(
  output        io_in_0_ready,
  input         io_in_0_valid,
  input         io_in_0_bits_threadId,
  input  [63:0] io_in_0_bits_programCounterOffset,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input         io_in_1_bits_threadId,
  input  [63:0] io_in_1_bits_programCounterOffset,
  input         io_out_ready,
  output        io_out_valid,
  output        io_out_bits_threadId,
  output [63:0] io_out_bits_programCounterOffset
);
  wire  grant_1 = ~io_in_0_valid; // @[Arbiter.scala 45:78]
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 146:19]
  assign io_in_1_ready = grant_1 & io_out_ready; // @[Arbiter.scala 146:19]
  assign io_out_valid = ~grant_1 | io_in_1_valid; // @[Arbiter.scala 147:31]
  assign io_out_bits_threadId = io_in_0_valid ? io_in_0_bits_threadId : io_in_1_bits_threadId; // @[Arbiter.scala 136:15 138:26 140:19]
  assign io_out_bits_programCounterOffset = io_in_0_valid ? $signed(io_in_0_bits_programCounterOffset) : $signed(
    io_in_1_bits_programCounterOffset); // @[Arbiter.scala 136:15 138:26 140:19]
endmodule
module BranchOutputCollector(
  input         clock,
  input         reset,
  output        io_fetch_0_addresses_valid,
  output        io_fetch_0_addresses_bits_threadId,
  output [63:0] io_fetch_0_addresses_bits_programCounterOffset,
  output        io_fetch_1_addresses_valid,
  output        io_fetch_1_addresses_bits_threadId,
  output [63:0] io_fetch_1_addresses_bits_programCounterOffset,
  output        io_executor_0_ready,
  input         io_executor_0_valid,
  input         io_executor_0_bits_threadId,
  input  [63:0] io_executor_0_bits_programCounterOffset,
  output        io_executor_1_ready,
  input         io_executor_1_valid,
  input         io_executor_1_bits_threadId,
  input  [63:0] io_executor_1_bits_programCounterOffset,
  input         io_isError_0,
  input         io_isError_1
);
  wire  threadFifos_0_clock; // @[BranchOutputCollector.scala 16:36]
  wire  threadFifos_0_reset; // @[BranchOutputCollector.scala 16:36]
  wire  threadFifos_0_input_ready; // @[BranchOutputCollector.scala 16:36]
  wire  threadFifos_0_input_valid; // @[BranchOutputCollector.scala 16:36]
  wire  threadFifos_0_input_bits_threadId; // @[BranchOutputCollector.scala 16:36]
  wire [63:0] threadFifos_0_input_bits_programCounterOffset; // @[BranchOutputCollector.scala 16:36]
  wire  threadFifos_0_output_valid; // @[BranchOutputCollector.scala 16:36]
  wire  threadFifos_0_output_bits_threadId; // @[BranchOutputCollector.scala 16:36]
  wire [63:0] threadFifos_0_output_bits_programCounterOffset; // @[BranchOutputCollector.scala 16:36]
  wire  threadFifos_0_flush; // @[BranchOutputCollector.scala 16:36]
  wire  threadFifos_1_clock; // @[BranchOutputCollector.scala 16:36]
  wire  threadFifos_1_reset; // @[BranchOutputCollector.scala 16:36]
  wire  threadFifos_1_input_ready; // @[BranchOutputCollector.scala 16:36]
  wire  threadFifos_1_input_valid; // @[BranchOutputCollector.scala 16:36]
  wire  threadFifos_1_input_bits_threadId; // @[BranchOutputCollector.scala 16:36]
  wire [63:0] threadFifos_1_input_bits_programCounterOffset; // @[BranchOutputCollector.scala 16:36]
  wire  threadFifos_1_output_valid; // @[BranchOutputCollector.scala 16:36]
  wire  threadFifos_1_output_bits_threadId; // @[BranchOutputCollector.scala 16:36]
  wire [63:0] threadFifos_1_output_bits_programCounterOffset; // @[BranchOutputCollector.scala 16:36]
  wire  threadFifos_1_flush; // @[BranchOutputCollector.scala 16:36]
  wire  executorArbiters_0_io_in_0_ready; // @[BranchOutputCollector.scala 18:11]
  wire  executorArbiters_0_io_in_0_valid; // @[BranchOutputCollector.scala 18:11]
  wire  executorArbiters_0_io_in_0_bits_threadId; // @[BranchOutputCollector.scala 18:11]
  wire [63:0] executorArbiters_0_io_in_0_bits_programCounterOffset; // @[BranchOutputCollector.scala 18:11]
  wire  executorArbiters_0_io_in_1_ready; // @[BranchOutputCollector.scala 18:11]
  wire  executorArbiters_0_io_in_1_valid; // @[BranchOutputCollector.scala 18:11]
  wire  executorArbiters_0_io_in_1_bits_threadId; // @[BranchOutputCollector.scala 18:11]
  wire [63:0] executorArbiters_0_io_in_1_bits_programCounterOffset; // @[BranchOutputCollector.scala 18:11]
  wire  executorArbiters_0_io_out_ready; // @[BranchOutputCollector.scala 18:11]
  wire  executorArbiters_0_io_out_valid; // @[BranchOutputCollector.scala 18:11]
  wire  executorArbiters_0_io_out_bits_threadId; // @[BranchOutputCollector.scala 18:11]
  wire [63:0] executorArbiters_0_io_out_bits_programCounterOffset; // @[BranchOutputCollector.scala 18:11]
  wire  executorArbiters_1_io_in_0_ready; // @[BranchOutputCollector.scala 18:11]
  wire  executorArbiters_1_io_in_0_valid; // @[BranchOutputCollector.scala 18:11]
  wire  executorArbiters_1_io_in_0_bits_threadId; // @[BranchOutputCollector.scala 18:11]
  wire [63:0] executorArbiters_1_io_in_0_bits_programCounterOffset; // @[BranchOutputCollector.scala 18:11]
  wire  executorArbiters_1_io_in_1_ready; // @[BranchOutputCollector.scala 18:11]
  wire  executorArbiters_1_io_in_1_valid; // @[BranchOutputCollector.scala 18:11]
  wire  executorArbiters_1_io_in_1_bits_threadId; // @[BranchOutputCollector.scala 18:11]
  wire [63:0] executorArbiters_1_io_in_1_bits_programCounterOffset; // @[BranchOutputCollector.scala 18:11]
  wire  executorArbiters_1_io_out_ready; // @[BranchOutputCollector.scala 18:11]
  wire  executorArbiters_1_io_out_valid; // @[BranchOutputCollector.scala 18:11]
  wire  executorArbiters_1_io_out_bits_threadId; // @[BranchOutputCollector.scala 18:11]
  wire [63:0] executorArbiters_1_io_out_bits_programCounterOffset; // @[BranchOutputCollector.scala 18:11]
  wire  _executorArbiters_0_io_in_0_valid_T = ~io_executor_0_bits_threadId; // @[BranchOutputCollector.scala 24:62]
  wire  _executorArbiters_0_io_in_1_valid_T = ~io_executor_1_bits_threadId; // @[BranchOutputCollector.scala 24:62]
  wire  _io_executor_0_ready_T_1 = executorArbiters_0_io_in_0_ready & _executorArbiters_0_io_in_0_valid_T; // @[BranchOutputCollector.scala 33:18]
  wire  _io_executor_0_ready_T_3 = executorArbiters_1_io_in_0_ready & io_executor_0_bits_threadId; // @[BranchOutputCollector.scala 33:18]
  wire  _io_executor_1_ready_T_1 = executorArbiters_0_io_in_1_ready & _executorArbiters_0_io_in_1_valid_T; // @[BranchOutputCollector.scala 33:18]
  wire  _io_executor_1_ready_T_3 = executorArbiters_1_io_in_1_ready & io_executor_1_bits_threadId; // @[BranchOutputCollector.scala 33:18]
  FIFO_3 threadFifos_0 ( // @[BranchOutputCollector.scala 16:36]
    .clock(threadFifos_0_clock),
    .reset(threadFifos_0_reset),
    .input_ready(threadFifos_0_input_ready),
    .input_valid(threadFifos_0_input_valid),
    .input_bits_threadId(threadFifos_0_input_bits_threadId),
    .input_bits_programCounterOffset(threadFifos_0_input_bits_programCounterOffset),
    .output_valid(threadFifos_0_output_valid),
    .output_bits_threadId(threadFifos_0_output_bits_threadId),
    .output_bits_programCounterOffset(threadFifos_0_output_bits_programCounterOffset),
    .flush(threadFifos_0_flush)
  );
  FIFO_3 threadFifos_1 ( // @[BranchOutputCollector.scala 16:36]
    .clock(threadFifos_1_clock),
    .reset(threadFifos_1_reset),
    .input_ready(threadFifos_1_input_ready),
    .input_valid(threadFifos_1_input_valid),
    .input_bits_threadId(threadFifos_1_input_bits_threadId),
    .input_bits_programCounterOffset(threadFifos_1_input_bits_programCounterOffset),
    .output_valid(threadFifos_1_output_valid),
    .output_bits_threadId(threadFifos_1_output_bits_threadId),
    .output_bits_programCounterOffset(threadFifos_1_output_bits_programCounterOffset),
    .flush(threadFifos_1_flush)
  );
  Arbiter_2 executorArbiters_0 ( // @[BranchOutputCollector.scala 18:11]
    .io_in_0_ready(executorArbiters_0_io_in_0_ready),
    .io_in_0_valid(executorArbiters_0_io_in_0_valid),
    .io_in_0_bits_threadId(executorArbiters_0_io_in_0_bits_threadId),
    .io_in_0_bits_programCounterOffset(executorArbiters_0_io_in_0_bits_programCounterOffset),
    .io_in_1_ready(executorArbiters_0_io_in_1_ready),
    .io_in_1_valid(executorArbiters_0_io_in_1_valid),
    .io_in_1_bits_threadId(executorArbiters_0_io_in_1_bits_threadId),
    .io_in_1_bits_programCounterOffset(executorArbiters_0_io_in_1_bits_programCounterOffset),
    .io_out_ready(executorArbiters_0_io_out_ready),
    .io_out_valid(executorArbiters_0_io_out_valid),
    .io_out_bits_threadId(executorArbiters_0_io_out_bits_threadId),
    .io_out_bits_programCounterOffset(executorArbiters_0_io_out_bits_programCounterOffset)
  );
  Arbiter_2 executorArbiters_1 ( // @[BranchOutputCollector.scala 18:11]
    .io_in_0_ready(executorArbiters_1_io_in_0_ready),
    .io_in_0_valid(executorArbiters_1_io_in_0_valid),
    .io_in_0_bits_threadId(executorArbiters_1_io_in_0_bits_threadId),
    .io_in_0_bits_programCounterOffset(executorArbiters_1_io_in_0_bits_programCounterOffset),
    .io_in_1_ready(executorArbiters_1_io_in_1_ready),
    .io_in_1_valid(executorArbiters_1_io_in_1_valid),
    .io_in_1_bits_threadId(executorArbiters_1_io_in_1_bits_threadId),
    .io_in_1_bits_programCounterOffset(executorArbiters_1_io_in_1_bits_programCounterOffset),
    .io_out_ready(executorArbiters_1_io_out_ready),
    .io_out_valid(executorArbiters_1_io_out_valid),
    .io_out_bits_threadId(executorArbiters_1_io_out_bits_threadId),
    .io_out_bits_programCounterOffset(executorArbiters_1_io_out_bits_programCounterOffset)
  );
  assign io_fetch_0_addresses_valid = threadFifos_0_output_valid; // @[BranchOutputCollector.scala 42:35]
  assign io_fetch_0_addresses_bits_threadId = threadFifos_0_output_bits_threadId; // @[BranchOutputCollector.scala 41:34]
  assign io_fetch_0_addresses_bits_programCounterOffset = threadFifos_0_output_bits_programCounterOffset; // @[BranchOutputCollector.scala 41:34]
  assign io_fetch_1_addresses_valid = threadFifos_1_output_valid; // @[BranchOutputCollector.scala 42:35]
  assign io_fetch_1_addresses_bits_threadId = threadFifos_1_output_bits_threadId; // @[BranchOutputCollector.scala 41:34]
  assign io_fetch_1_addresses_bits_programCounterOffset = threadFifos_1_output_bits_programCounterOffset; // @[BranchOutputCollector.scala 41:34]
  assign io_executor_0_ready = _io_executor_0_ready_T_1 | _io_executor_0_ready_T_3; // @[BranchOutputCollector.scala 35:17]
  assign io_executor_1_ready = _io_executor_1_ready_T_1 | _io_executor_1_ready_T_3; // @[BranchOutputCollector.scala 35:17]
  assign threadFifos_0_clock = clock;
  assign threadFifos_0_reset = reset;
  assign threadFifos_0_input_valid = executorArbiters_0_io_out_valid; // @[BranchOutputCollector.scala 39:28]
  assign threadFifos_0_input_bits_threadId = executorArbiters_0_io_out_bits_threadId; // @[BranchOutputCollector.scala 39:28]
  assign threadFifos_0_input_bits_programCounterOffset = executorArbiters_0_io_out_bits_programCounterOffset; // @[BranchOutputCollector.scala 39:28]
  assign threadFifos_0_flush = io_isError_0; // @[BranchOutputCollector.scala 40:28]
  assign threadFifos_1_clock = clock;
  assign threadFifos_1_reset = reset;
  assign threadFifos_1_input_valid = executorArbiters_1_io_out_valid; // @[BranchOutputCollector.scala 39:28]
  assign threadFifos_1_input_bits_threadId = executorArbiters_1_io_out_bits_threadId; // @[BranchOutputCollector.scala 39:28]
  assign threadFifos_1_input_bits_programCounterOffset = executorArbiters_1_io_out_bits_programCounterOffset; // @[BranchOutputCollector.scala 39:28]
  assign threadFifos_1_flush = io_isError_1; // @[BranchOutputCollector.scala 40:28]
  assign executorArbiters_0_io_in_0_valid = io_executor_0_valid & ~io_executor_0_bits_threadId; // @[BranchOutputCollector.scala 24:30]
  assign executorArbiters_0_io_in_0_bits_threadId = io_executor_0_bits_threadId; // @[BranchOutputCollector.scala 22:38]
  assign executorArbiters_0_io_in_0_bits_programCounterOffset = io_executor_0_bits_programCounterOffset; // @[BranchOutputCollector.scala 22:38]
  assign executorArbiters_0_io_in_1_valid = io_executor_1_valid & ~io_executor_1_bits_threadId; // @[BranchOutputCollector.scala 24:30]
  assign executorArbiters_0_io_in_1_bits_threadId = io_executor_1_bits_threadId; // @[BranchOutputCollector.scala 22:38]
  assign executorArbiters_0_io_in_1_bits_programCounterOffset = io_executor_1_bits_programCounterOffset; // @[BranchOutputCollector.scala 22:38]
  assign executorArbiters_0_io_out_ready = threadFifos_0_input_ready; // @[BranchOutputCollector.scala 39:28]
  assign executorArbiters_1_io_in_0_valid = io_executor_0_valid & io_executor_0_bits_threadId; // @[BranchOutputCollector.scala 24:30]
  assign executorArbiters_1_io_in_0_bits_threadId = io_executor_0_bits_threadId; // @[BranchOutputCollector.scala 22:38]
  assign executorArbiters_1_io_in_0_bits_programCounterOffset = io_executor_0_bits_programCounterOffset; // @[BranchOutputCollector.scala 22:38]
  assign executorArbiters_1_io_in_1_valid = io_executor_1_valid & io_executor_1_bits_threadId; // @[BranchOutputCollector.scala 24:30]
  assign executorArbiters_1_io_in_1_bits_threadId = io_executor_1_bits_threadId; // @[BranchOutputCollector.scala 22:38]
  assign executorArbiters_1_io_in_1_bits_programCounterOffset = io_executor_1_bits_programCounterOffset; // @[BranchOutputCollector.scala 22:38]
  assign executorArbiters_1_io_out_ready = threadFifos_1_input_ready; // @[BranchOutputCollector.scala 39:28]
endmodule
module Uncompresser(
  output        io_fetch_ready,
  input         io_fetch_valid,
  input  [31:0] io_fetch_bits_instruction,
  input  [63:0] io_fetch_bits_programCounter,
  input         io_decoder_ready,
  output        io_decoder_valid,
  output [31:0] io_decoder_bits_instruction,
  output [63:0] io_decoder_bits_programCounter,
  output        io_decoder_bits_wasCompressed
);
  wire  _io_decoder_bits_instruction_T_3 = io_fetch_bits_instruction[12:2] != 11'h0; // @[Uncompresser.scala 188:32]
  wire [9:0] _io_decoder_bits_instruction_T_10 = {io_fetch_bits_instruction[10:7],io_fetch_bits_instruction[12:11],
    io_fetch_bits_instruction[5],io_fetch_bits_instruction[6],2'h0}; // @[Cat.scala 33:92]
  wire [11:0] io_decoder_bits_instruction_w = {{2'd0}, _io_decoder_bits_instruction_T_10}; // @[Uncompresser.scala 160:17 161:7]
  wire [31:0] io_decoder_bits_instruction_output = {io_decoder_bits_instruction_w,5'h2,3'h0,2'h1,
    io_fetch_bits_instruction[4:2],7'h13}; // @[Uncompresser.scala 19:51]
  wire [31:0] _io_decoder_bits_instruction_T_11 = _io_decoder_bits_instruction_T_3 ? io_decoder_bits_instruction_output
     : 32'h0; // @[Uncompresser.scala 187:26]
  wire [6:0] _io_decoder_bits_instruction_T_19 = {io_fetch_bits_instruction[5],io_fetch_bits_instruction[12:10],
    io_fetch_bits_instruction[6],2'h0}; // @[Cat.scala 33:92]
  wire [11:0] io_decoder_bits_instruction_w_1 = {{5'd0}, _io_decoder_bits_instruction_T_19}; // @[Uncompresser.scala 160:17 161:7]
  wire [31:0] io_decoder_bits_instruction_output_1 = {io_decoder_bits_instruction_w_1,2'h1,io_fetch_bits_instruction[9:7
    ],3'h2,2'h1,io_fetch_bits_instruction[4:2],7'h3}; // @[Uncompresser.scala 19:51]
  wire [7:0] _io_decoder_bits_instruction_T_26 = {io_fetch_bits_instruction[6:5],io_fetch_bits_instruction[12:10],3'h0}; // @[Cat.scala 33:92]
  wire [11:0] io_decoder_bits_instruction_w_2 = {{4'd0}, _io_decoder_bits_instruction_T_26}; // @[Uncompresser.scala 160:17 161:7]
  wire [31:0] io_decoder_bits_instruction_output_2 = {io_decoder_bits_instruction_w_2,2'h1,io_fetch_bits_instruction[9:7
    ],3'h3,2'h1,io_fetch_bits_instruction[4:2],7'h3}; // @[Uncompresser.scala 19:51]
  wire [31:0] io_decoder_bits_instruction_output_3 = {io_decoder_bits_instruction_w_1[11:5],2'h1,
    io_fetch_bits_instruction[4:2],2'h1,io_fetch_bits_instruction[9:7],3'h2,io_decoder_bits_instruction_w_1[4:0],7'h23}; // @[Uncompresser.scala 60:61]
  wire [31:0] io_decoder_bits_instruction_output_4 = {io_decoder_bits_instruction_w_2[11:5],2'h1,
    io_fetch_bits_instruction[4:2],2'h1,io_fetch_bits_instruction[9:7],3'h3,io_decoder_bits_instruction_w_2[4:0],7'h23}; // @[Uncompresser.scala 60:61]
  wire [31:0] _io_decoder_bits_instruction_T_43 = 3'h0 == io_fetch_bits_instruction[15:13] ?
    _io_decoder_bits_instruction_T_11 : 32'h0; // @[Mux.scala 81:58]
  wire [31:0] _io_decoder_bits_instruction_T_45 = 3'h2 == io_fetch_bits_instruction[15:13] ?
    io_decoder_bits_instruction_output_1 : _io_decoder_bits_instruction_T_43; // @[Mux.scala 81:58]
  wire [31:0] _io_decoder_bits_instruction_T_47 = 3'h3 == io_fetch_bits_instruction[15:13] ?
    io_decoder_bits_instruction_output_2 : _io_decoder_bits_instruction_T_45; // @[Mux.scala 81:58]
  wire [31:0] _io_decoder_bits_instruction_T_49 = 3'h6 == io_fetch_bits_instruction[15:13] ?
    io_decoder_bits_instruction_output_3 : _io_decoder_bits_instruction_T_47; // @[Mux.scala 81:58]
  wire [31:0] _io_decoder_bits_instruction_T_51 = 3'h7 == io_fetch_bits_instruction[15:13] ?
    io_decoder_bits_instruction_output_4 : _io_decoder_bits_instruction_T_49; // @[Mux.scala 81:58]
  wire  _io_decoder_bits_instruction_T_54 = io_fetch_bits_instruction[11:7] == 5'h0; // @[Uncompresser.scala 259:32]
  wire [5:0] _io_decoder_bits_instruction_T_59 = {io_fetch_bits_instruction[12],io_fetch_bits_instruction[6:2]}; // @[Uncompresser.scala 265:42]
  wire  _io_decoder_bits_instruction_w_T_1 = ~_io_decoder_bits_instruction_T_59[5]; // @[Uncompresser.scala 150:7]
  wire [11:0] _io_decoder_bits_instruction_w_T_3 = {6'h3f,io_fetch_bits_instruction[12],io_fetch_bits_instruction[6:2]}; // @[Uncompresser.scala 152:39]
  wire [11:0] io_decoder_bits_instruction_w_5 = _io_decoder_bits_instruction_w_T_1 ? {{6'd0},
    _io_decoder_bits_instruction_T_59} : _io_decoder_bits_instruction_w_T_3; // @[Uncompresser.scala 149:13]
  wire [31:0] io_decoder_bits_instruction_output_6 = {io_decoder_bits_instruction_w_5,io_fetch_bits_instruction[11:7],3'h0
    ,io_fetch_bits_instruction[11:7],7'h13}; // @[Uncompresser.scala 19:51]
  wire [31:0] _io_decoder_bits_instruction_T_60 = _io_decoder_bits_instruction_T_54 ? 32'h13 :
    io_decoder_bits_instruction_output_6; // @[Uncompresser.scala 258:26]
  wire [31:0] io_decoder_bits_instruction_output_7 = {io_decoder_bits_instruction_w_5,io_fetch_bits_instruction[11:7],3'h0
    ,io_fetch_bits_instruction[11:7],7'h1b}; // @[Uncompresser.scala 19:51]
  wire [31:0] _io_decoder_bits_instruction_T_68 = _io_decoder_bits_instruction_T_54 ? 32'h0 :
    io_decoder_bits_instruction_output_7; // @[Uncompresser.scala 268:26]
  wire [31:0] io_decoder_bits_instruction_output_8 = {io_decoder_bits_instruction_w_5,5'h0,3'h0,
    io_fetch_bits_instruction[11:7],7'h13}; // @[Uncompresser.scala 19:51]
  wire [31:0] _io_decoder_bits_instruction_T_75 = _io_decoder_bits_instruction_T_54 ? 32'h0 :
    io_decoder_bits_instruction_output_8; // @[Uncompresser.scala 278:26]
  wire  _io_decoder_bits_instruction_T_77 = io_fetch_bits_instruction[11:7] == 5'h2; // @[Uncompresser.scala 291:35]
  wire [9:0] _io_decoder_bits_instruction_T_83 = {io_fetch_bits_instruction[12],io_fetch_bits_instruction[4:3],
    io_fetch_bits_instruction[5],io_fetch_bits_instruction[2],io_fetch_bits_instruction[6],4'h0}; // @[Cat.scala 33:92]
  wire  _io_decoder_bits_instruction_w_T_16 = ~_io_decoder_bits_instruction_T_83[9]; // @[Uncompresser.scala 150:7]
  wire [11:0] _io_decoder_bits_instruction_w_T_18 = {2'h3,io_fetch_bits_instruction[12],io_fetch_bits_instruction[4:3],
    io_fetch_bits_instruction[5],io_fetch_bits_instruction[2],io_fetch_bits_instruction[6],4'h0}; // @[Uncompresser.scala 152:39]
  wire [11:0] io_decoder_bits_instruction_w_8 = _io_decoder_bits_instruction_w_T_16 ? {{2'd0},
    _io_decoder_bits_instruction_T_83} : _io_decoder_bits_instruction_w_T_18; // @[Uncompresser.scala 149:13]
  wire [31:0] io_decoder_bits_instruction_output_9 = {io_decoder_bits_instruction_w_8,5'h2,3'h0,5'h2,7'h13}; // @[Uncompresser.scala 19:51]
  wire  _io_decoder_bits_instruction_T_85 = io_fetch_bits_instruction[11:7] != 5'h2; // @[Uncompresser.scala 307:35]
  wire [19:0] _io_decoder_bits_instruction_w_T_23 = {14'h3fff,io_fetch_bits_instruction[12],io_fetch_bits_instruction[6:
    2]}; // @[Uncompresser.scala 152:39]
  wire [19:0] io_decoder_bits_instruction_w_9 = _io_decoder_bits_instruction_w_T_1 ? {{14'd0},
    _io_decoder_bits_instruction_T_59} : _io_decoder_bits_instruction_w_T_23; // @[Uncompresser.scala 149:13]
  wire [31:0] io_decoder_bits_instruction_output_10 = {io_decoder_bits_instruction_w_9,io_fetch_bits_instruction[11:7],7'h37
    }; // @[Uncompresser.scala 110:28]
  wire [31:0] _io_decoder_bits_instruction_T_90 = _io_decoder_bits_instruction_T_85 ?
    io_decoder_bits_instruction_output_10 : 32'h0; // @[Mux.scala 101:16]
  wire [31:0] _io_decoder_bits_instruction_T_91 = _io_decoder_bits_instruction_T_77 ?
    io_decoder_bits_instruction_output_9 : _io_decoder_bits_instruction_T_90; // @[Mux.scala 101:16]
  wire [31:0] io_decoder_bits_instruction_output_11 = {6'h0,io_fetch_bits_instruction[12],io_fetch_bits_instruction[6:2]
    ,2'h1,io_fetch_bits_instruction[9:7],3'h5,2'h1,io_fetch_bits_instruction[9:7],7'h13}; // @[Uncompresser.scala 37:56]
  wire [31:0] io_decoder_bits_instruction_output_12 = {6'h10,io_fetch_bits_instruction[12],io_fetch_bits_instruction[6:2
    ],2'h1,io_fetch_bits_instruction[9:7],3'h5,2'h1,io_fetch_bits_instruction[9:7],7'h13}; // @[Uncompresser.scala 37:56]
  wire [31:0] io_decoder_bits_instruction_output_13 = {io_decoder_bits_instruction_w_5,2'h1,io_fetch_bits_instruction[9:
    7],3'h7,2'h1,io_fetch_bits_instruction[9:7],7'h13}; // @[Uncompresser.scala 19:51]
  wire [31:0] io_decoder_bits_instruction_output_14 = {7'h20,2'h1,io_fetch_bits_instruction[4:2],2'h1,
    io_fetch_bits_instruction[9:7],3'h0,2'h1,io_fetch_bits_instruction[9:7],7'h3b}; // @[Uncompresser.scala 132:56]
  wire [31:0] io_decoder_bits_instruction_output_15 = {7'h0,2'h1,io_fetch_bits_instruction[4:2],2'h1,
    io_fetch_bits_instruction[9:7],3'h0,2'h1,io_fetch_bits_instruction[9:7],7'h3b}; // @[Uncompresser.scala 132:56]
  wire [31:0] _io_decoder_bits_instruction_T_129 = 2'h0 == io_fetch_bits_instruction[6:5] ?
    io_decoder_bits_instruction_output_14 : 32'h0; // @[Mux.scala 81:58]
  wire [31:0] _io_decoder_bits_instruction_T_131 = 2'h1 == io_fetch_bits_instruction[6:5] ?
    io_decoder_bits_instruction_output_15 : _io_decoder_bits_instruction_T_129; // @[Mux.scala 81:58]
  wire [31:0] io_decoder_bits_instruction_output_16 = {7'h20,2'h1,io_fetch_bits_instruction[4:2],2'h1,
    io_fetch_bits_instruction[9:7],3'h0,2'h1,io_fetch_bits_instruction[9:7],7'h33}; // @[Uncompresser.scala 132:56]
  wire [31:0] io_decoder_bits_instruction_output_17 = {7'h0,2'h1,io_fetch_bits_instruction[4:2],2'h1,
    io_fetch_bits_instruction[9:7],3'h4,2'h1,io_fetch_bits_instruction[9:7],7'h33}; // @[Uncompresser.scala 132:56]
  wire [31:0] io_decoder_bits_instruction_output_18 = {7'h0,2'h1,io_fetch_bits_instruction[4:2],2'h1,
    io_fetch_bits_instruction[9:7],3'h6,2'h1,io_fetch_bits_instruction[9:7],7'h33}; // @[Uncompresser.scala 132:56]
  wire [31:0] io_decoder_bits_instruction_output_19 = {7'h0,2'h1,io_fetch_bits_instruction[4:2],2'h1,
    io_fetch_bits_instruction[9:7],3'h7,2'h1,io_fetch_bits_instruction[9:7],7'h33}; // @[Uncompresser.scala 132:56]
  wire [31:0] _io_decoder_bits_instruction_T_158 = 2'h1 == io_fetch_bits_instruction[6:5] ?
    io_decoder_bits_instruction_output_17 : io_decoder_bits_instruction_output_16; // @[Mux.scala 81:58]
  wire [31:0] _io_decoder_bits_instruction_T_160 = 2'h2 == io_fetch_bits_instruction[6:5] ?
    io_decoder_bits_instruction_output_18 : _io_decoder_bits_instruction_T_158; // @[Mux.scala 81:58]
  wire [31:0] _io_decoder_bits_instruction_T_162 = 2'h3 == io_fetch_bits_instruction[6:5] ?
    io_decoder_bits_instruction_output_19 : _io_decoder_bits_instruction_T_160; // @[Mux.scala 81:58]
  wire [31:0] _io_decoder_bits_instruction_T_163 = io_fetch_bits_instruction[12] ? _io_decoder_bits_instruction_T_131 :
    _io_decoder_bits_instruction_T_162; // @[Uncompresser.scala 336:29]
  wire [31:0] _io_decoder_bits_instruction_T_165 = 2'h1 == io_fetch_bits_instruction[11:10] ?
    io_decoder_bits_instruction_output_12 : io_decoder_bits_instruction_output_11; // @[Mux.scala 81:58]
  wire [31:0] _io_decoder_bits_instruction_T_167 = 2'h2 == io_fetch_bits_instruction[11:10] ?
    io_decoder_bits_instruction_output_13 : _io_decoder_bits_instruction_T_165; // @[Mux.scala 81:58]
  wire [31:0] _io_decoder_bits_instruction_T_169 = 2'h3 == io_fetch_bits_instruction[11:10] ?
    _io_decoder_bits_instruction_T_163 : _io_decoder_bits_instruction_T_167; // @[Mux.scala 81:58]
  wire [11:0] _io_decoder_bits_instruction_T_178 = {io_fetch_bits_instruction[12],io_fetch_bits_instruction[8],
    io_fetch_bits_instruction[10:9],io_fetch_bits_instruction[6],io_fetch_bits_instruction[7],io_fetch_bits_instruction[
    2],io_fetch_bits_instruction[11],io_fetch_bits_instruction[5:3],1'h0}; // @[Cat.scala 33:92]
  wire  _io_decoder_bits_instruction_w_T_31 = ~_io_decoder_bits_instruction_T_178[11]; // @[Uncompresser.scala 150:7]
  wire [21:0] _io_decoder_bits_instruction_w_T_33 = {10'h3ff,io_fetch_bits_instruction[12],io_fetch_bits_instruction[8],
    io_fetch_bits_instruction[10:9],io_fetch_bits_instruction[6],io_fetch_bits_instruction[7],io_fetch_bits_instruction[
    2],io_fetch_bits_instruction[11],io_fetch_bits_instruction[5:3],1'h0}; // @[Uncompresser.scala 152:39]
  wire [21:0] io_decoder_bits_instruction_w_13 = _io_decoder_bits_instruction_w_T_31 ? {{10'd0},
    _io_decoder_bits_instruction_T_178} : _io_decoder_bits_instruction_w_T_33; // @[Uncompresser.scala 149:13]
  wire [31:0] io_decoder_bits_instruction_output_20 = {io_decoder_bits_instruction_w_13[20],
    io_decoder_bits_instruction_w_13[10:1],io_decoder_bits_instruction_w_13[11],io_decoder_bits_instruction_w_13[19:12],5'h0
    ,7'h6f}; // @[Cat.scala 33:92]
  wire [8:0] _io_decoder_bits_instruction_T_186 = {io_fetch_bits_instruction[12],io_fetch_bits_instruction[6:5],
    io_fetch_bits_instruction[2],io_fetch_bits_instruction[11:10],io_fetch_bits_instruction[4:3],1'h0}; // @[Cat.scala 33:92]
  wire  _io_decoder_bits_instruction_w_T_36 = ~_io_decoder_bits_instruction_T_186[8]; // @[Uncompresser.scala 150:7]
  wire [12:0] _io_decoder_bits_instruction_w_T_38 = {4'hf,io_fetch_bits_instruction[12],io_fetch_bits_instruction[6:5],
    io_fetch_bits_instruction[2],io_fetch_bits_instruction[11:10],io_fetch_bits_instruction[4:3],1'h0}; // @[Uncompresser.scala 152:39]
  wire [12:0] io_decoder_bits_instruction_w_14 = _io_decoder_bits_instruction_w_T_36 ? {{4'd0},
    _io_decoder_bits_instruction_T_186} : _io_decoder_bits_instruction_w_T_38; // @[Uncompresser.scala 149:13]
  wire [31:0] io_decoder_bits_instruction_output_21 = {io_decoder_bits_instruction_w_14[12],
    io_decoder_bits_instruction_w_14[10:5],5'h0,2'h1,io_fetch_bits_instruction[9:7],3'h0,
    io_decoder_bits_instruction_w_14[4:1],io_decoder_bits_instruction_w_14[11],7'h63}; // @[Uncompresser.scala 83:18]
  wire [31:0] io_decoder_bits_instruction_output_22 = {io_decoder_bits_instruction_w_14[12],
    io_decoder_bits_instruction_w_14[10:5],5'h0,2'h1,io_fetch_bits_instruction[9:7],3'h1,
    io_decoder_bits_instruction_w_14[4:1],io_decoder_bits_instruction_w_14[11],7'h63}; // @[Uncompresser.scala 83:18]
  wire [31:0] _io_decoder_bits_instruction_T_196 = 3'h1 == io_fetch_bits_instruction[15:13] ?
    _io_decoder_bits_instruction_T_68 : _io_decoder_bits_instruction_T_60; // @[Mux.scala 81:58]
  wire [31:0] _io_decoder_bits_instruction_T_198 = 3'h2 == io_fetch_bits_instruction[15:13] ?
    _io_decoder_bits_instruction_T_75 : _io_decoder_bits_instruction_T_196; // @[Mux.scala 81:58]
  wire [31:0] _io_decoder_bits_instruction_T_200 = 3'h3 == io_fetch_bits_instruction[15:13] ?
    _io_decoder_bits_instruction_T_91 : _io_decoder_bits_instruction_T_198; // @[Mux.scala 81:58]
  wire [31:0] _io_decoder_bits_instruction_T_202 = 3'h4 == io_fetch_bits_instruction[15:13] ?
    _io_decoder_bits_instruction_T_169 : _io_decoder_bits_instruction_T_200; // @[Mux.scala 81:58]
  wire [31:0] _io_decoder_bits_instruction_T_204 = 3'h5 == io_fetch_bits_instruction[15:13] ?
    io_decoder_bits_instruction_output_20 : _io_decoder_bits_instruction_T_202; // @[Mux.scala 81:58]
  wire [31:0] _io_decoder_bits_instruction_T_206 = 3'h6 == io_fetch_bits_instruction[15:13] ?
    io_decoder_bits_instruction_output_21 : _io_decoder_bits_instruction_T_204; // @[Mux.scala 81:58]
  wire [31:0] _io_decoder_bits_instruction_T_208 = 3'h7 == io_fetch_bits_instruction[15:13] ?
    io_decoder_bits_instruction_output_22 : _io_decoder_bits_instruction_T_206; // @[Mux.scala 81:58]
  wire [31:0] io_decoder_bits_instruction_output_23 = {6'h0,io_fetch_bits_instruction[12],io_fetch_bits_instruction[6:2]
    ,io_fetch_bits_instruction[11:7],3'h1,io_fetch_bits_instruction[11:7],7'h13}; // @[Uncompresser.scala 37:56]
  wire [7:0] _io_decoder_bits_instruction_T_219 = {io_fetch_bits_instruction[3:2],io_fetch_bits_instruction[12],
    io_fetch_bits_instruction[6:4],2'h0}; // @[Cat.scala 33:92]
  wire [11:0] io_decoder_bits_instruction_w_17 = {{4'd0}, _io_decoder_bits_instruction_T_219}; // @[Uncompresser.scala 160:17 161:7]
  wire [31:0] io_decoder_bits_instruction_output_24 = {io_decoder_bits_instruction_w_17,5'h2,3'h2,
    io_fetch_bits_instruction[11:7],7'h3}; // @[Uncompresser.scala 19:51]
  wire [8:0] _io_decoder_bits_instruction_T_224 = {io_fetch_bits_instruction[4:2],io_fetch_bits_instruction[12],
    io_fetch_bits_instruction[6:5],3'h0}; // @[Cat.scala 33:92]
  wire [11:0] io_decoder_bits_instruction_w_18 = {{3'd0}, _io_decoder_bits_instruction_T_224}; // @[Uncompresser.scala 160:17 161:7]
  wire [31:0] io_decoder_bits_instruction_output_25 = {io_decoder_bits_instruction_w_18,5'h2,3'h3,
    io_fetch_bits_instruction[11:7],7'h3}; // @[Uncompresser.scala 19:51]
  wire  _io_decoder_bits_instruction_T_226 = ~io_fetch_bits_instruction[12]; // @[Uncompresser.scala 480:13]
  wire  _io_decoder_bits_instruction_T_228 = io_fetch_bits_instruction[6:2] == 5'h0; // @[Uncompresser.scala 482:33]
  wire [31:0] io_decoder_bits_instruction_output_26 = {12'h0,io_fetch_bits_instruction[11:7],3'h0,5'h0,7'h67}; // @[Uncompresser.scala 19:51]
  wire [31:0] io_decoder_bits_instruction_output_27 = {12'h0,io_fetch_bits_instruction[6:2],3'h0,
    io_fetch_bits_instruction[11:7],7'h13}; // @[Uncompresser.scala 19:51]
  wire [31:0] _io_decoder_bits_instruction_T_232 = _io_decoder_bits_instruction_T_228 ?
    io_decoder_bits_instruction_output_26 : io_decoder_bits_instruction_output_27; // @[Uncompresser.scala 481:16]
  wire [31:0] io_decoder_bits_instruction_output_28 = {12'h0,io_fetch_bits_instruction[11:7],3'h0,5'h1,7'h67}; // @[Uncompresser.scala 19:51]
  wire [31:0] io_decoder_bits_instruction_output_29 = {7'h0,io_fetch_bits_instruction[6:2],io_fetch_bits_instruction[11:
    7],3'h0,io_fetch_bits_instruction[11:7],7'h33}; // @[Uncompresser.scala 132:56]
  wire [31:0] _io_decoder_bits_instruction_T_241 = _io_decoder_bits_instruction_T_228 ?
    io_decoder_bits_instruction_output_28 : io_decoder_bits_instruction_output_29; // @[Uncompresser.scala 494:18]
  wire [31:0] _io_decoder_bits_instruction_T_242 = _io_decoder_bits_instruction_T_54 ? 32'h0 :
    _io_decoder_bits_instruction_T_241; // @[Uncompresser.scala 491:16]
  wire [31:0] _io_decoder_bits_instruction_T_243 = _io_decoder_bits_instruction_T_226 ?
    _io_decoder_bits_instruction_T_232 : _io_decoder_bits_instruction_T_242; // @[Uncompresser.scala 479:26]
  wire [7:0] _io_decoder_bits_instruction_T_247 = {io_fetch_bits_instruction[8:7],io_fetch_bits_instruction[12:9],2'h0}; // @[Cat.scala 33:92]
  wire [11:0] io_decoder_bits_instruction_w_19 = {{4'd0}, _io_decoder_bits_instruction_T_247}; // @[Uncompresser.scala 160:17 161:7]
  wire [31:0] io_decoder_bits_instruction_output_30 = {io_decoder_bits_instruction_w_19[11:5],io_fetch_bits_instruction[
    6:2],5'h2,3'h2,io_decoder_bits_instruction_w_19[4:0],7'h23}; // @[Uncompresser.scala 60:61]
  wire [8:0] _io_decoder_bits_instruction_T_251 = {io_fetch_bits_instruction[9:7],io_fetch_bits_instruction[12:10],3'h0}
    ; // @[Cat.scala 33:92]
  wire [11:0] io_decoder_bits_instruction_w_20 = {{3'd0}, _io_decoder_bits_instruction_T_251}; // @[Uncompresser.scala 160:17 161:7]
  wire [31:0] io_decoder_bits_instruction_output_31 = {io_decoder_bits_instruction_w_20[11:5],io_fetch_bits_instruction[
    6:2],5'h2,3'h3,io_decoder_bits_instruction_w_20[4:0],7'h23}; // @[Uncompresser.scala 60:61]
  wire [31:0] _io_decoder_bits_instruction_T_253 = 3'h0 == io_fetch_bits_instruction[15:13] ?
    io_decoder_bits_instruction_output_23 : 32'h0; // @[Mux.scala 81:58]
  wire [31:0] _io_decoder_bits_instruction_T_255 = 3'h2 == io_fetch_bits_instruction[15:13] ?
    io_decoder_bits_instruction_output_24 : _io_decoder_bits_instruction_T_253; // @[Mux.scala 81:58]
  wire [31:0] _io_decoder_bits_instruction_T_257 = 3'h3 == io_fetch_bits_instruction[15:13] ?
    io_decoder_bits_instruction_output_25 : _io_decoder_bits_instruction_T_255; // @[Mux.scala 81:58]
  wire [31:0] _io_decoder_bits_instruction_T_259 = 3'h4 == io_fetch_bits_instruction[15:13] ?
    _io_decoder_bits_instruction_T_243 : _io_decoder_bits_instruction_T_257; // @[Mux.scala 81:58]
  wire [31:0] _io_decoder_bits_instruction_T_261 = 3'h6 == io_fetch_bits_instruction[15:13] ?
    io_decoder_bits_instruction_output_30 : _io_decoder_bits_instruction_T_259; // @[Mux.scala 81:58]
  wire [31:0] _io_decoder_bits_instruction_T_263 = 3'h7 == io_fetch_bits_instruction[15:13] ?
    io_decoder_bits_instruction_output_31 : _io_decoder_bits_instruction_T_261; // @[Mux.scala 81:58]
  wire [31:0] _io_decoder_bits_instruction_T_265 = 2'h1 == io_fetch_bits_instruction[1:0] ?
    _io_decoder_bits_instruction_T_208 : _io_decoder_bits_instruction_T_51; // @[Mux.scala 81:58]
  wire [31:0] _io_decoder_bits_instruction_T_267 = 2'h2 == io_fetch_bits_instruction[1:0] ?
    _io_decoder_bits_instruction_T_263 : _io_decoder_bits_instruction_T_265; // @[Mux.scala 81:58]
  assign io_fetch_ready = io_decoder_ready; // @[Uncompresser.scala 172:18]
  assign io_decoder_valid = io_fetch_valid; // @[Uncompresser.scala 173:20]
  assign io_decoder_bits_instruction = 2'h3 == io_fetch_bits_instruction[1:0] ? io_fetch_bits_instruction :
    _io_decoder_bits_instruction_T_267; // @[Mux.scala 81:58]
  assign io_decoder_bits_programCounter = io_fetch_bits_programCounter; // @[Uncompresser.scala 174:34]
  assign io_decoder_bits_wasCompressed = io_fetch_bits_instruction[1:0] != 2'h3; // @[Uncompresser.scala 178:54]
endmodule
module OpcodeFormatChecker(
  input  [6:0] io_opcode,
  output [2:0] io_format
);
  wire [2:0] _io_format_T_1 = 7'h3 == io_opcode ? 3'h1 : 3'h6; // @[Mux.scala 81:58]
  wire [2:0] _io_format_T_3 = 7'hf == io_opcode ? 3'h1 : _io_format_T_1; // @[Mux.scala 81:58]
  wire [2:0] _io_format_T_5 = 7'h73 == io_opcode ? 3'h1 : _io_format_T_3; // @[Mux.scala 81:58]
  wire [2:0] _io_format_T_7 = 7'h13 == io_opcode ? 3'h1 : _io_format_T_5; // @[Mux.scala 81:58]
  wire [2:0] _io_format_T_9 = 7'h1b == io_opcode ? 3'h1 : _io_format_T_7; // @[Mux.scala 81:58]
  wire [2:0] _io_format_T_11 = 7'h67 == io_opcode ? 3'h1 : _io_format_T_9; // @[Mux.scala 81:58]
  wire [2:0] _io_format_T_13 = 7'h6f == io_opcode ? 3'h2 : _io_format_T_11; // @[Mux.scala 81:58]
  wire [2:0] _io_format_T_15 = 7'h37 == io_opcode ? 3'h4 : _io_format_T_13; // @[Mux.scala 81:58]
  wire [2:0] _io_format_T_17 = 7'h17 == io_opcode ? 3'h4 : _io_format_T_15; // @[Mux.scala 81:58]
  wire [2:0] _io_format_T_19 = 7'h63 == io_opcode ? 3'h5 : _io_format_T_17; // @[Mux.scala 81:58]
  wire [2:0] _io_format_T_21 = 7'h23 == io_opcode ? 3'h3 : _io_format_T_19; // @[Mux.scala 81:58]
  wire [2:0] _io_format_T_23 = 7'h33 == io_opcode ? 3'h0 : _io_format_T_21; // @[Mux.scala 81:58]
  assign io_format = 7'h3b == io_opcode ? 3'h0 : _io_format_T_23; // @[Mux.scala 81:58]
endmodule
module SourceTagSelector(
  input        io_reorderBufferDestinationTag_valid,
  input        io_reorderBufferDestinationTag_bits_threadId,
  input  [3:0] io_reorderBufferDestinationTag_bits_id,
  output       io_sourceTag_valid,
  output       io_sourceTag_tag_threadId,
  output [3:0] io_sourceTag_tag_id
);
  assign io_sourceTag_valid = io_reorderBufferDestinationTag_valid; // @[SourceTagSelector.scala 35:56]
  assign io_sourceTag_tag_threadId = io_sourceTag_valid & io_reorderBufferDestinationTag_bits_threadId; // @[SourceTagSelector.scala 43:28 44:22 60:22]
  assign io_sourceTag_tag_id = io_sourceTag_valid ? io_reorderBufferDestinationTag_bits_id : 4'h0; // @[SourceTagSelector.scala 43:28 44:22 60:22]
endmodule
module ValueSelector1(
  input         io_reorderBufferValue_valid,
  input  [63:0] io_reorderBufferValue_bits,
  input  [63:0] io_registerFileValue,
  input         io_outputCollector_outputs_valid,
  input         io_outputCollector_outputs_bits_resultType,
  input  [63:0] io_outputCollector_outputs_bits_value,
  input         io_outputCollector_outputs_bits_tag_threadId,
  input  [3:0]  io_outputCollector_outputs_bits_tag_id,
  input  [63:0] io_immediateValue,
  input  [2:0]  io_opcodeFormat,
  input         io_sourceTag_valid,
  input         io_sourceTag_tag_threadId,
  input  [3:0]  io_sourceTag_tag_id,
  output        io_value_valid,
  output [63:0] io_value_bits
);
  wire  _outputMatchingTagExists_T_4 = io_outputCollector_outputs_bits_tag_id == io_sourceTag_tag_id &
    io_outputCollector_outputs_bits_tag_threadId == io_sourceTag_tag_threadId; // @[Tag.scala 13:25]
  wire  outputMatchingTagExists = io_outputCollector_outputs_valid & ~io_outputCollector_outputs_bits_resultType &
    _outputMatchingTagExists_T_4; // @[ValueSelector1.scala 29:56]
  wire  _io_value_valid_T = io_opcodeFormat == 3'h4; // @[ValueSelector1.scala 35:24]
  wire  _io_value_valid_T_1 = io_opcodeFormat == 3'h2; // @[ValueSelector1.scala 35:49]
  wire  _io_value_valid_T_2 = io_opcodeFormat == 3'h4 | io_opcodeFormat == 3'h2; // @[ValueSelector1.scala 35:30]
  wire  _io_value_valid_T_4 = io_sourceTag_valid & io_reorderBufferValue_valid; // @[ValueSelector1.scala 37:27]
  wire  _io_value_valid_T_5 = io_sourceTag_valid & outputMatchingTagExists; // @[ValueSelector1.scala 38:27]
  wire  _io_value_valid_T_6 = ~io_sourceTag_valid; // @[ValueSelector1.scala 39:8]
  wire [63:0] _io_value_bits_T_8 = _io_value_valid_T_6 ? io_registerFileValue : 64'h0; // @[Mux.scala 101:16]
  wire [63:0] _io_value_bits_T_9 = _io_value_valid_T_5 ? io_outputCollector_outputs_bits_value : _io_value_bits_T_8; // @[Mux.scala 101:16]
  wire [63:0] _io_value_bits_T_10 = _io_value_valid_T_4 ? io_reorderBufferValue_bits : _io_value_bits_T_9; // @[Mux.scala 101:16]
  wire [63:0] _io_value_bits_T_12 = _io_value_valid_T_1 ? io_immediateValue : _io_value_bits_T_10; // @[Mux.scala 101:16]
  assign io_value_valid = _io_value_valid_T_2 | (_io_value_valid_T_4 | (_io_value_valid_T_5 | _io_value_valid_T_6)); // @[Mux.scala 101:16]
  assign io_value_bits = _io_value_valid_T ? io_immediateValue : _io_value_bits_T_12; // @[Mux.scala 101:16]
endmodule
module ValueSelector2(
  input         io_reorderBufferValue_valid,
  input  [63:0] io_reorderBufferValue_bits,
  input  [63:0] io_registerFileValue,
  input  [63:0] io_programCounter,
  input         io_outputCollector_outputs_valid,
  input         io_outputCollector_outputs_bits_resultType,
  input  [63:0] io_outputCollector_outputs_bits_value,
  input         io_outputCollector_outputs_bits_tag_threadId,
  input  [3:0]  io_outputCollector_outputs_bits_tag_id,
  input  [2:0]  io_opcodeFormat,
  input         io_sourceTag_valid,
  input         io_sourceTag_tag_threadId,
  input  [3:0]  io_sourceTag_tag_id,
  output        io_value_valid,
  output [63:0] io_value_bits
);
  wire  _outputMatchingTagExists_T_4 = io_outputCollector_outputs_bits_tag_id == io_sourceTag_tag_id &
    io_outputCollector_outputs_bits_tag_threadId == io_sourceTag_tag_threadId; // @[Tag.scala 13:25]
  wire  outputMatchingTagExists = io_outputCollector_outputs_valid & ~io_outputCollector_outputs_bits_resultType &
    _outputMatchingTagExists_T_4; // @[ValueSelector2.scala 28:56]
  wire  _io_value_valid_T = io_opcodeFormat == 3'h1; // @[ValueSelector2.scala 34:24]
  wire  _io_value_valid_T_1 = io_opcodeFormat == 3'h4; // @[ValueSelector2.scala 34:49]
  wire  _io_value_valid_T_3 = io_opcodeFormat == 3'h2; // @[ValueSelector2.scala 34:74]
  wire  _io_value_valid_T_4 = io_opcodeFormat == 3'h1 | io_opcodeFormat == 3'h4 | io_opcodeFormat == 3'h2; // @[ValueSelector2.scala 34:55]
  wire  _io_value_valid_T_6 = io_sourceTag_valid & io_reorderBufferValue_valid; // @[ValueSelector2.scala 36:27]
  wire  _io_value_valid_T_7 = io_sourceTag_valid & outputMatchingTagExists; // @[ValueSelector2.scala 37:27]
  wire  _io_value_valid_T_8 = ~io_sourceTag_valid; // @[ValueSelector2.scala 38:8]
  wire  _io_value_bits_T_4 = _io_value_valid_T | _io_value_valid_T_3 | _io_value_valid_T_1; // @[ValueSelector2.scala 44:55]
  wire [63:0] _io_value_bits_T_9 = _io_value_valid_T_8 ? io_registerFileValue : 64'h0; // @[Mux.scala 101:16]
  wire [63:0] _io_value_bits_T_10 = _io_value_valid_T_7 ? io_outputCollector_outputs_bits_value : _io_value_bits_T_9; // @[Mux.scala 101:16]
  wire [63:0] _io_value_bits_T_11 = _io_value_valid_T_6 ? io_reorderBufferValue_bits : _io_value_bits_T_10; // @[Mux.scala 101:16]
  assign io_value_valid = _io_value_valid_T_4 | (_io_value_valid_T_6 | (_io_value_valid_T_7 | _io_value_valid_T_8)); // @[Mux.scala 101:16]
  assign io_value_bits = _io_value_bits_T_4 ? io_programCounter : _io_value_bits_T_11; // @[Mux.scala 101:16]
endmodule
module Decoder(
  output        io_instructionFetch_ready,
  input         io_instructionFetch_valid,
  input  [31:0] io_instructionFetch_bits_instruction,
  input  [63:0] io_instructionFetch_bits_programCounter,
  input         io_instructionFetch_bits_wasCompressed,
  output [4:0]  io_reorderBuffer_source1_sourceRegister,
  input         io_reorderBuffer_source1_matchingTag_valid,
  input  [3:0]  io_reorderBuffer_source1_matchingTag_bits_id,
  input         io_reorderBuffer_source1_value_valid,
  input  [63:0] io_reorderBuffer_source1_value_bits,
  output [4:0]  io_reorderBuffer_source2_sourceRegister,
  input         io_reorderBuffer_source2_matchingTag_valid,
  input  [3:0]  io_reorderBuffer_source2_matchingTag_bits_id,
  input         io_reorderBuffer_source2_value_valid,
  input  [63:0] io_reorderBuffer_source2_value_bits,
  output [4:0]  io_reorderBuffer_destination_destinationRegister,
  input  [3:0]  io_reorderBuffer_destination_destinationTag_id,
  output        io_reorderBuffer_destination_storeSign,
  input         io_reorderBuffer_ready,
  output        io_reorderBuffer_valid,
  input         io_outputCollector_outputs_valid,
  input         io_outputCollector_outputs_bits_resultType,
  input  [63:0] io_outputCollector_outputs_bits_value,
  input         io_outputCollector_outputs_bits_tag_threadId,
  input  [3:0]  io_outputCollector_outputs_bits_tag_id,
  output [4:0]  io_registerFile_sourceRegister1,
  output [4:0]  io_registerFile_sourceRegister2,
  input  [63:0] io_registerFile_value1,
  input  [63:0] io_registerFile_value2,
  input         io_reservationStation_ready,
  output [6:0]  io_reservationStation_entry_opcode,
  output [2:0]  io_reservationStation_entry_function3,
  output [11:0] io_reservationStation_entry_immediateOrFunction7,
  output        io_reservationStation_entry_sourceTag1_threadId,
  output [3:0]  io_reservationStation_entry_sourceTag1_id,
  output        io_reservationStation_entry_ready1,
  output [63:0] io_reservationStation_entry_value1,
  output        io_reservationStation_entry_sourceTag2_threadId,
  output [3:0]  io_reservationStation_entry_sourceTag2_id,
  output        io_reservationStation_entry_ready2,
  output [63:0] io_reservationStation_entry_value2,
  output        io_reservationStation_entry_destinationTag_threadId,
  output [3:0]  io_reservationStation_entry_destinationTag_id,
  output        io_reservationStation_entry_wasCompressed,
  output        io_reservationStation_entry_valid,
  input         io_loadStoreQueue_ready,
  output        io_loadStoreQueue_valid,
  output        io_loadStoreQueue_bits_accessInfo_accessType,
  output        io_loadStoreQueue_bits_accessInfo_signed,
  output [1:0]  io_loadStoreQueue_bits_accessInfo_accessWidth,
  output        io_loadStoreQueue_bits_addressAndLoadResultTag_threadId,
  output [3:0]  io_loadStoreQueue_bits_addressAndLoadResultTag_id,
  output [63:0] io_loadStoreQueue_bits_address,
  output        io_loadStoreQueue_bits_addressValid,
  output        io_loadStoreQueue_bits_storeDataTag_threadId,
  output [3:0]  io_loadStoreQueue_bits_storeDataTag_id,
  output [63:0] io_loadStoreQueue_bits_storeData,
  output        io_loadStoreQueue_bits_storeDataValid,
  input         io_csr_ready,
  output        io_csr_valid,
  output        io_csr_bits_sourceTag_threadId,
  output [3:0]  io_csr_bits_sourceTag_id,
  output [3:0]  io_csr_bits_destinationTag_id,
  output [63:0] io_csr_bits_value,
  output        io_csr_bits_ready,
  output [11:0] io_csr_bits_address,
  output [1:0]  io_csr_bits_csrAccessType
);
  wire [6:0] opcodeFormatChecker_io_opcode; // @[Decoder.scala 78:35]
  wire [2:0] opcodeFormatChecker_io_format; // @[Decoder.scala 78:35]
  wire  sourceTagSelector1_io_reorderBufferDestinationTag_valid; // @[Decoder.scala 126:34]
  wire  sourceTagSelector1_io_reorderBufferDestinationTag_bits_threadId; // @[Decoder.scala 126:34]
  wire [3:0] sourceTagSelector1_io_reorderBufferDestinationTag_bits_id; // @[Decoder.scala 126:34]
  wire  sourceTagSelector1_io_sourceTag_valid; // @[Decoder.scala 126:34]
  wire  sourceTagSelector1_io_sourceTag_tag_threadId; // @[Decoder.scala 126:34]
  wire [3:0] sourceTagSelector1_io_sourceTag_tag_id; // @[Decoder.scala 126:34]
  wire  sourceTagSelector2_io_reorderBufferDestinationTag_valid; // @[Decoder.scala 141:34]
  wire  sourceTagSelector2_io_reorderBufferDestinationTag_bits_threadId; // @[Decoder.scala 141:34]
  wire [3:0] sourceTagSelector2_io_reorderBufferDestinationTag_bits_id; // @[Decoder.scala 141:34]
  wire  sourceTagSelector2_io_sourceTag_valid; // @[Decoder.scala 141:34]
  wire  sourceTagSelector2_io_sourceTag_tag_threadId; // @[Decoder.scala 141:34]
  wire [3:0] sourceTagSelector2_io_sourceTag_tag_id; // @[Decoder.scala 141:34]
  wire  valueSelector1_io_reorderBufferValue_valid; // @[Decoder.scala 155:30]
  wire [63:0] valueSelector1_io_reorderBufferValue_bits; // @[Decoder.scala 155:30]
  wire [63:0] valueSelector1_io_registerFileValue; // @[Decoder.scala 155:30]
  wire  valueSelector1_io_outputCollector_outputs_valid; // @[Decoder.scala 155:30]
  wire  valueSelector1_io_outputCollector_outputs_bits_resultType; // @[Decoder.scala 155:30]
  wire [63:0] valueSelector1_io_outputCollector_outputs_bits_value; // @[Decoder.scala 155:30]
  wire  valueSelector1_io_outputCollector_outputs_bits_tag_threadId; // @[Decoder.scala 155:30]
  wire [3:0] valueSelector1_io_outputCollector_outputs_bits_tag_id; // @[Decoder.scala 155:30]
  wire [63:0] valueSelector1_io_immediateValue; // @[Decoder.scala 155:30]
  wire [2:0] valueSelector1_io_opcodeFormat; // @[Decoder.scala 155:30]
  wire  valueSelector1_io_sourceTag_valid; // @[Decoder.scala 155:30]
  wire  valueSelector1_io_sourceTag_tag_threadId; // @[Decoder.scala 155:30]
  wire [3:0] valueSelector1_io_sourceTag_tag_id; // @[Decoder.scala 155:30]
  wire  valueSelector1_io_value_valid; // @[Decoder.scala 155:30]
  wire [63:0] valueSelector1_io_value_bits; // @[Decoder.scala 155:30]
  wire  valueSelector2_io_reorderBufferValue_valid; // @[Decoder.scala 167:30]
  wire [63:0] valueSelector2_io_reorderBufferValue_bits; // @[Decoder.scala 167:30]
  wire [63:0] valueSelector2_io_registerFileValue; // @[Decoder.scala 167:30]
  wire [63:0] valueSelector2_io_programCounter; // @[Decoder.scala 167:30]
  wire  valueSelector2_io_outputCollector_outputs_valid; // @[Decoder.scala 167:30]
  wire  valueSelector2_io_outputCollector_outputs_bits_resultType; // @[Decoder.scala 167:30]
  wire [63:0] valueSelector2_io_outputCollector_outputs_bits_value; // @[Decoder.scala 167:30]
  wire  valueSelector2_io_outputCollector_outputs_bits_tag_threadId; // @[Decoder.scala 167:30]
  wire [3:0] valueSelector2_io_outputCollector_outputs_bits_tag_id; // @[Decoder.scala 167:30]
  wire [2:0] valueSelector2_io_opcodeFormat; // @[Decoder.scala 167:30]
  wire  valueSelector2_io_sourceTag_valid; // @[Decoder.scala 167:30]
  wire  valueSelector2_io_sourceTag_tag_threadId; // @[Decoder.scala 167:30]
  wire [3:0] valueSelector2_io_sourceTag_tag_id; // @[Decoder.scala 167:30]
  wire  valueSelector2_io_value_valid; // @[Decoder.scala 167:30]
  wire [63:0] valueSelector2_io_value_bits; // @[Decoder.scala 167:30]
  wire [4:0] instRd = io_instructionFetch_bits_instruction[11:7]; // @[Decoder.scala 46:52]
  wire [4:0] instRs1 = io_instructionFetch_bits_instruction[19:15]; // @[Decoder.scala 47:53]
  wire [4:0] instRs2 = io_instructionFetch_bits_instruction[24:20]; // @[Decoder.scala 48:53]
  wire [2:0] instFunct3 = io_instructionFetch_bits_instruction[14:12]; // @[Decoder.scala 49:56]
  wire [6:0] instFunct7 = io_instructionFetch_bits_instruction[31:25]; // @[Decoder.scala 50:56]
  wire [6:0] instOp = io_instructionFetch_bits_instruction[6:0]; // @[Decoder.scala 51:52]
  wire [11:0] instImmS = {instFunct7,instRd}; // @[Cat.scala 33:92]
  wire [11:0] instImmB = {io_instructionFetch_bits_instruction[31],io_instructionFetch_bits_instruction[7],
    io_instructionFetch_bits_instruction[30:25],io_instructionFetch_bits_instruction[11:8]}; // @[Cat.scala 33:92]
  wire [19:0] instImmU = io_instructionFetch_bits_instruction[31:12]; // @[Decoder.scala 63:54]
  wire [11:0] immIExtended = io_instructionFetch_bits_instruction[31:20]; // @[Decoder.scala 73:14]
  wire [31:0] immUExtended = {instImmU,12'h0}; // @[Decoder.scala 74:47]
  wire [20:0] immJExtended = {io_instructionFetch_bits_instruction[31],io_instructionFetch_bits_instruction[19:12],
    io_instructionFetch_bits_instruction[20],io_instructionFetch_bits_instruction[30:21],1'h0}; // @[Decoder.scala 75:46]
  wire  _destinationIsValid_T = opcodeFormatChecker_io_format == 3'h0; // @[Decoder.scala 82:58]
  wire  _destinationIsValid_T_1 = opcodeFormatChecker_io_format == 3'h1; // @[Decoder.scala 83:35]
  wire  _destinationIsValid_T_2 = opcodeFormatChecker_io_format == 3'h0 | _destinationIsValid_T_1; // @[Decoder.scala 82:64]
  wire  _destinationIsValid_T_3 = opcodeFormatChecker_io_format == 3'h4; // @[Decoder.scala 84:35]
  wire  _destinationIsValid_T_4 = _destinationIsValid_T_2 | _destinationIsValid_T_3; // @[Decoder.scala 83:41]
  wire  _destinationIsValid_T_5 = opcodeFormatChecker_io_format == 3'h2; // @[Decoder.scala 85:35]
  wire  destinationIsValid = _destinationIsValid_T_4 | _destinationIsValid_T_5; // @[Decoder.scala 84:41]
  wire  _source1IsValid_T_3 = opcodeFormatChecker_io_format == 3'h3; // @[Decoder.scala 90:35]
  wire  _source1IsValid_T_4 = _destinationIsValid_T_2 | _source1IsValid_T_3; // @[Decoder.scala 89:41]
  wire  _source1IsValid_T_5 = opcodeFormatChecker_io_format == 3'h5; // @[Decoder.scala 91:35]
  wire  source1IsValid = _source1IsValid_T_4 | _source1IsValid_T_5; // @[Decoder.scala 90:41]
  wire  _source2IsValid_T_2 = _destinationIsValid_T | _source1IsValid_T_3; // @[Decoder.scala 94:60]
  wire  source2IsValid = _source2IsValid_T_2 | _source1IsValid_T_5; // @[Decoder.scala 95:41]
  wire  _io_reorderBuffer_destination_storeSign_T = instOp == 7'h23; // @[Decoder.scala 106:52]
  wire [2:0] _valueSelector1_io_immediateValue_T = opcodeFormatChecker_io_format; // @[Decoder.scala 162:35]
  wire [31:0] _valueSelector1_io_immediateValue_T_4 = 3'h4 == _valueSelector1_io_immediateValue_T ? $signed(immUExtended
    ) : $signed(32'sh0); // @[Mux.scala 81:58]
  wire [31:0] _valueSelector1_io_immediateValue_T_6 = 3'h2 == _valueSelector1_io_immediateValue_T ? $signed({{11{
    immJExtended[20]}},immJExtended}) : $signed(_valueSelector1_io_immediateValue_T_4); // @[Mux.scala 81:58]
  wire  _io_reorderBuffer_valid_T = io_instructionFetch_ready & io_instructionFetch_valid; // @[Decoder.scala 194:55]
  wire [6:0] _io_reservationStation_entry_valid_T_1 = instOp & 7'h5f; // @[Decoder.scala 197:14]
  wire  _io_reservationStation_entry_valid_T_2 = 7'h3 == _io_reservationStation_entry_valid_T_1; // @[Decoder.scala 197:14]
  wire  _io_reservationStation_entry_valid_T_3 = _io_reservationStation_entry_valid_T_2 & valueSelector1_io_value_valid; // @[Decoder.scala 199:7]
  wire  _io_reservationStation_entry_valid_T_4 = ~_io_reservationStation_entry_valid_T_3; // @[Decoder.scala 197:5]
  wire  _io_reservationStation_entry_valid_T_5 = _io_reorderBuffer_valid_T & _io_reservationStation_entry_valid_T_4; // @[Decoder.scala 196:31]
  wire [11:0] _io_reservationStation_entry_immediateOrFunction7_T_2 = {instFunct7,5'h0}; // @[Cat.scala 33:92]
  wire [11:0] _io_reservationStation_entry_immediateOrFunction7_T_6 = io_instructionFetch_bits_instruction[31:20]; // @[Decoder.scala 212:32]
  wire [11:0] _io_reservationStation_entry_immediateOrFunction7_T_8 = 3'h0 == _valueSelector1_io_immediateValue_T ?
    _io_reservationStation_entry_immediateOrFunction7_T_2 : 12'h0; // @[Mux.scala 81:58]
  wire [11:0] _io_reservationStation_entry_immediateOrFunction7_T_10 = 3'h3 == _valueSelector1_io_immediateValue_T ?
    instImmS : _io_reservationStation_entry_immediateOrFunction7_T_8; // @[Mux.scala 81:58]
  wire [11:0] _io_reservationStation_entry_immediateOrFunction7_T_12 = 3'h5 == _valueSelector1_io_immediateValue_T ?
    instImmB : _io_reservationStation_entry_immediateOrFunction7_T_10; // @[Mux.scala 81:58]
  wire  _io_loadStoreQueue_valid_T_2 = io_loadStoreQueue_ready & _io_reservationStation_entry_valid_T_2; // @[Decoder.scala 233:54]
  wire  _io_loadStoreQueue_bits_accessInfo_w_accessWidth_T_3 = instFunct3[1:0] == 2'h1; // @[MemoryAccessWidth.scala 13:23]
  wire  _io_loadStoreQueue_bits_accessInfo_w_accessWidth_T_5 = instFunct3[1:0] == 2'h2; // @[MemoryAccessWidth.scala 14:23]
  wire  _io_loadStoreQueue_bits_accessInfo_w_accessWidth_T_7 = instFunct3[1:0] == 2'h3; // @[MemoryAccessWidth.scala 15:23]
  wire [1:0] _io_loadStoreQueue_bits_accessInfo_w_accessWidth_T_13 =
    _io_loadStoreQueue_bits_accessInfo_w_accessWidth_T_5 ? 2'h2 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_loadStoreQueue_bits_accessInfo_w_accessWidth_T_15 =
    _io_loadStoreQueue_bits_accessInfo_w_accessWidth_T_7 ? 2'h3 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _GEN_27 = {{1'd0}, _io_loadStoreQueue_bits_accessInfo_w_accessWidth_T_3}; // @[Mux.scala 27:73]
  wire [1:0] _io_loadStoreQueue_bits_accessInfo_w_accessWidth_T_17 = _GEN_27 |
    _io_loadStoreQueue_bits_accessInfo_w_accessWidth_T_13; // @[Mux.scala 27:73]
  wire [11:0] _io_loadStoreQueue_bits_address_T_2 = {instFunct7,instRd}; // @[Decoder.scala 245:16]
  wire [11:0] _io_loadStoreQueue_bits_address_T_4 = _io_reorderBuffer_destination_storeSign_T ? $signed(
    _io_loadStoreQueue_bits_address_T_2) : $signed(immIExtended); // @[Decoder.scala 243:81]
  wire [63:0] _GEN_28 = {{52{_io_loadStoreQueue_bits_address_T_4[11]}},_io_loadStoreQueue_bits_address_T_4}; // @[Decoder.scala 243:76]
  OpcodeFormatChecker opcodeFormatChecker ( // @[Decoder.scala 78:35]
    .io_opcode(opcodeFormatChecker_io_opcode),
    .io_format(opcodeFormatChecker_io_format)
  );
  SourceTagSelector sourceTagSelector1 ( // @[Decoder.scala 126:34]
    .io_reorderBufferDestinationTag_valid(sourceTagSelector1_io_reorderBufferDestinationTag_valid),
    .io_reorderBufferDestinationTag_bits_threadId(sourceTagSelector1_io_reorderBufferDestinationTag_bits_threadId),
    .io_reorderBufferDestinationTag_bits_id(sourceTagSelector1_io_reorderBufferDestinationTag_bits_id),
    .io_sourceTag_valid(sourceTagSelector1_io_sourceTag_valid),
    .io_sourceTag_tag_threadId(sourceTagSelector1_io_sourceTag_tag_threadId),
    .io_sourceTag_tag_id(sourceTagSelector1_io_sourceTag_tag_id)
  );
  SourceTagSelector sourceTagSelector2 ( // @[Decoder.scala 141:34]
    .io_reorderBufferDestinationTag_valid(sourceTagSelector2_io_reorderBufferDestinationTag_valid),
    .io_reorderBufferDestinationTag_bits_threadId(sourceTagSelector2_io_reorderBufferDestinationTag_bits_threadId),
    .io_reorderBufferDestinationTag_bits_id(sourceTagSelector2_io_reorderBufferDestinationTag_bits_id),
    .io_sourceTag_valid(sourceTagSelector2_io_sourceTag_valid),
    .io_sourceTag_tag_threadId(sourceTagSelector2_io_sourceTag_tag_threadId),
    .io_sourceTag_tag_id(sourceTagSelector2_io_sourceTag_tag_id)
  );
  ValueSelector1 valueSelector1 ( // @[Decoder.scala 155:30]
    .io_reorderBufferValue_valid(valueSelector1_io_reorderBufferValue_valid),
    .io_reorderBufferValue_bits(valueSelector1_io_reorderBufferValue_bits),
    .io_registerFileValue(valueSelector1_io_registerFileValue),
    .io_outputCollector_outputs_valid(valueSelector1_io_outputCollector_outputs_valid),
    .io_outputCollector_outputs_bits_resultType(valueSelector1_io_outputCollector_outputs_bits_resultType),
    .io_outputCollector_outputs_bits_value(valueSelector1_io_outputCollector_outputs_bits_value),
    .io_outputCollector_outputs_bits_tag_threadId(valueSelector1_io_outputCollector_outputs_bits_tag_threadId),
    .io_outputCollector_outputs_bits_tag_id(valueSelector1_io_outputCollector_outputs_bits_tag_id),
    .io_immediateValue(valueSelector1_io_immediateValue),
    .io_opcodeFormat(valueSelector1_io_opcodeFormat),
    .io_sourceTag_valid(valueSelector1_io_sourceTag_valid),
    .io_sourceTag_tag_threadId(valueSelector1_io_sourceTag_tag_threadId),
    .io_sourceTag_tag_id(valueSelector1_io_sourceTag_tag_id),
    .io_value_valid(valueSelector1_io_value_valid),
    .io_value_bits(valueSelector1_io_value_bits)
  );
  ValueSelector2 valueSelector2 ( // @[Decoder.scala 167:30]
    .io_reorderBufferValue_valid(valueSelector2_io_reorderBufferValue_valid),
    .io_reorderBufferValue_bits(valueSelector2_io_reorderBufferValue_bits),
    .io_registerFileValue(valueSelector2_io_registerFileValue),
    .io_programCounter(valueSelector2_io_programCounter),
    .io_outputCollector_outputs_valid(valueSelector2_io_outputCollector_outputs_valid),
    .io_outputCollector_outputs_bits_resultType(valueSelector2_io_outputCollector_outputs_bits_resultType),
    .io_outputCollector_outputs_bits_value(valueSelector2_io_outputCollector_outputs_bits_value),
    .io_outputCollector_outputs_bits_tag_threadId(valueSelector2_io_outputCollector_outputs_bits_tag_threadId),
    .io_outputCollector_outputs_bits_tag_id(valueSelector2_io_outputCollector_outputs_bits_tag_id),
    .io_opcodeFormat(valueSelector2_io_opcodeFormat),
    .io_sourceTag_valid(valueSelector2_io_sourceTag_valid),
    .io_sourceTag_tag_threadId(valueSelector2_io_sourceTag_tag_threadId),
    .io_sourceTag_tag_id(valueSelector2_io_sourceTag_tag_id),
    .io_value_valid(valueSelector2_io_value_valid),
    .io_value_bits(valueSelector2_io_value_bits)
  );
  assign io_instructionFetch_ready = io_reservationStation_ready & io_reorderBuffer_ready & io_loadStoreQueue_ready &
    io_csr_ready; // @[Decoder.scala 192:113]
  assign io_reorderBuffer_source1_sourceRegister = source1IsValid ? instRs1 : 5'h0; // @[Decoder.scala 99:49]
  assign io_reorderBuffer_source2_sourceRegister = source2IsValid ? instRs2 : 5'h0; // @[Decoder.scala 100:49]
  assign io_reorderBuffer_destination_destinationRegister = destinationIsValid ? instRd : 5'h0; // @[Decoder.scala 101:58]
  assign io_reorderBuffer_destination_storeSign = instOp == 7'h23; // @[Decoder.scala 106:52]
  assign io_reorderBuffer_valid = io_instructionFetch_ready & io_instructionFetch_valid; // @[Decoder.scala 194:55]
  assign io_registerFile_sourceRegister1 = io_instructionFetch_bits_instruction[19:15]; // @[Decoder.scala 47:53]
  assign io_registerFile_sourceRegister2 = io_instructionFetch_bits_instruction[24:20]; // @[Decoder.scala 48:53]
  assign io_reservationStation_entry_opcode = io_instructionFetch_bits_instruction[6:0]; // @[Decoder.scala 51:52]
  assign io_reservationStation_entry_function3 = io_instructionFetch_bits_instruction[14:12]; // @[Decoder.scala 49:56]
  assign io_reservationStation_entry_immediateOrFunction7 = 3'h1 == _valueSelector1_io_immediateValue_T ?
    _io_reservationStation_entry_immediateOrFunction7_T_6 : _io_reservationStation_entry_immediateOrFunction7_T_12; // @[Mux.scala 81:58]
  assign io_reservationStation_entry_sourceTag1_threadId = valueSelector1_io_value_valid ? 1'h0 :
    sourceTagSelector1_io_sourceTag_tag_threadId; // @[Decoder.scala 216:23]
  assign io_reservationStation_entry_sourceTag1_id = valueSelector1_io_value_valid ? 4'h0 :
    sourceTagSelector1_io_sourceTag_tag_id; // @[Decoder.scala 216:23]
  assign io_reservationStation_entry_ready1 = valueSelector1_io_value_valid; // @[Decoder.scala 226:13]
  assign io_reservationStation_entry_value1 = valueSelector1_io_value_bits; // @[Decoder.scala 228:13]
  assign io_reservationStation_entry_sourceTag2_threadId = valueSelector2_io_value_valid ? 1'h0 :
    sourceTagSelector2_io_sourceTag_tag_threadId; // @[Decoder.scala 221:23]
  assign io_reservationStation_entry_sourceTag2_id = valueSelector2_io_value_valid ? 4'h0 :
    sourceTagSelector2_io_sourceTag_tag_id; // @[Decoder.scala 221:23]
  assign io_reservationStation_entry_ready2 = valueSelector2_io_value_valid; // @[Decoder.scala 227:13]
  assign io_reservationStation_entry_value2 = valueSelector2_io_value_bits; // @[Decoder.scala 229:13]
  assign io_reservationStation_entry_destinationTag_threadId = 1'h0; // @[Decoder.scala 215:21]
  assign io_reservationStation_entry_destinationTag_id = io_reorderBuffer_destination_destinationTag_id; // @[Decoder.scala 215:21]
  assign io_reservationStation_entry_wasCompressed = io_instructionFetch_bits_wasCompressed; // @[Decoder.scala 230:20]
  assign io_reservationStation_entry_valid = _io_reservationStation_entry_valid_T_5 & instOp != 7'h73; // @[Decoder.scala 199:41]
  assign io_loadStoreQueue_valid = _io_loadStoreQueue_valid_T_2 & io_instructionFetch_ready & io_instructionFetch_valid; // @[Decoder.scala 235:34]
  assign io_loadStoreQueue_bits_accessInfo_accessType = ~instOp[5]; // @[MemoryAccessType.scala 15:20]
  assign io_loadStoreQueue_bits_accessInfo_signed = ~instFunct3[2]; // @[MemoryAccessInfo.scala 15:17]
  assign io_loadStoreQueue_bits_accessInfo_accessWidth = _io_loadStoreQueue_bits_accessInfo_w_accessWidth_T_17 |
    _io_loadStoreQueue_bits_accessInfo_w_accessWidth_T_15; // @[Mux.scala 27:73]
  assign io_loadStoreQueue_bits_addressAndLoadResultTag_threadId = io_reservationStation_entry_destinationTag_threadId; // @[Decoder.scala 239:33 241:52]
  assign io_loadStoreQueue_bits_addressAndLoadResultTag_id = io_reservationStation_entry_destinationTag_id; // @[Decoder.scala 239:33 241:52]
  assign io_loadStoreQueue_bits_address = $signed(valueSelector1_io_value_bits) + $signed(_GEN_28); // @[Decoder.scala 247:8]
  assign io_loadStoreQueue_bits_addressValid = valueSelector1_io_value_valid; // @[Decoder.scala 239:33 242:41]
  assign io_loadStoreQueue_bits_storeDataTag_threadId = _io_reorderBuffer_destination_storeSign_T &
    valueSelector2_io_sourceTag_tag_threadId; // @[Decoder.scala 248:28 249:43 253:43]
  assign io_loadStoreQueue_bits_storeDataTag_id = _io_reorderBuffer_destination_storeSign_T ?
    valueSelector2_io_sourceTag_tag_id : 4'h0; // @[Decoder.scala 248:28 249:43 253:43]
  assign io_loadStoreQueue_bits_storeData = _io_reorderBuffer_destination_storeSign_T ? valueSelector2_io_value_bits : 64'h0
    ; // @[Decoder.scala 248:28 250:40 254:40]
  assign io_loadStoreQueue_bits_storeDataValid = _io_reorderBuffer_destination_storeSign_T ?
    valueSelector2_io_value_valid : 1'h1; // @[Decoder.scala 248:28 251:45 255:45]
  assign io_csr_valid = io_csr_ready & io_instructionFetch_ready & io_instructionFetch_valid & 7'h73 == instOp &
    instFunct3 != 3'h0; // @[Decoder.scala 261:117]
  assign io_csr_bits_sourceTag_threadId = valueSelector1_io_sourceTag_tag_threadId; // @[Decoder.scala 263:22 274:27]
  assign io_csr_bits_sourceTag_id = valueSelector1_io_sourceTag_tag_id; // @[Decoder.scala 263:22 274:27]
  assign io_csr_bits_destinationTag_id = io_reorderBuffer_destination_destinationTag_id; // @[Decoder.scala 263:22 285:32]
  assign io_csr_bits_value = instFunct3[2] ? {{59'd0}, instRs1} : valueSelector1_io_value_bits; // @[Decoder.scala 275:29]
  assign io_csr_bits_ready = instFunct3[2] | valueSelector1_io_value_valid; // @[Decoder.scala 280:29]
  assign io_csr_bits_address = io_instructionFetch_bits_instruction[31:20]; // @[Decoder.scala 52:54]
  assign io_csr_bits_csrAccessType = 2'h3 == instFunct3[1:0] ? 2'h2 : {{1'd0}, 2'h2 == instFunct3[1:0]}; // @[Mux.scala 81:58]
  assign opcodeFormatChecker_io_opcode = io_instructionFetch_bits_instruction[6:0]; // @[Decoder.scala 51:52]
  assign sourceTagSelector1_io_reorderBufferDestinationTag_valid = io_reorderBuffer_source1_matchingTag_valid; // @[Decoder.scala 127:53]
  assign sourceTagSelector1_io_reorderBufferDestinationTag_bits_threadId = 1'h0; // @[Decoder.scala 127:53]
  assign sourceTagSelector1_io_reorderBufferDestinationTag_bits_id = io_reorderBuffer_source1_matchingTag_bits_id; // @[Decoder.scala 127:53]
  assign sourceTagSelector2_io_reorderBufferDestinationTag_valid = io_reorderBuffer_source2_matchingTag_valid; // @[Decoder.scala 142:53]
  assign sourceTagSelector2_io_reorderBufferDestinationTag_bits_threadId = 1'h0; // @[Decoder.scala 142:53]
  assign sourceTagSelector2_io_reorderBufferDestinationTag_bits_id = io_reorderBuffer_source2_matchingTag_bits_id; // @[Decoder.scala 142:53]
  assign valueSelector1_io_reorderBufferValue_valid = io_reorderBuffer_source1_value_valid; // @[Decoder.scala 157:40]
  assign valueSelector1_io_reorderBufferValue_bits = io_reorderBuffer_source1_value_bits; // @[Decoder.scala 157:40]
  assign valueSelector1_io_registerFileValue = io_registerFile_value1; // @[Decoder.scala 158:39]
  assign valueSelector1_io_outputCollector_outputs_valid = io_outputCollector_outputs_valid; // @[Decoder.scala 159:37]
  assign valueSelector1_io_outputCollector_outputs_bits_resultType = io_outputCollector_outputs_bits_resultType; // @[Decoder.scala 159:37]
  assign valueSelector1_io_outputCollector_outputs_bits_value = io_outputCollector_outputs_bits_value; // @[Decoder.scala 159:37]
  assign valueSelector1_io_outputCollector_outputs_bits_tag_threadId = io_outputCollector_outputs_bits_tag_threadId; // @[Decoder.scala 159:37]
  assign valueSelector1_io_outputCollector_outputs_bits_tag_id = io_outputCollector_outputs_bits_tag_id; // @[Decoder.scala 159:37]
  assign valueSelector1_io_immediateValue = {{32{_valueSelector1_io_immediateValue_T_6[31]}},
    _valueSelector1_io_immediateValue_T_6}; // @[Decoder.scala 161:36]
  assign valueSelector1_io_opcodeFormat = opcodeFormatChecker_io_format; // @[Decoder.scala 160:34]
  assign valueSelector1_io_sourceTag_valid = sourceTagSelector1_io_sourceTag_valid; // @[Decoder.scala 156:31]
  assign valueSelector1_io_sourceTag_tag_threadId = sourceTagSelector1_io_sourceTag_tag_threadId; // @[Decoder.scala 156:31]
  assign valueSelector1_io_sourceTag_tag_id = sourceTagSelector1_io_sourceTag_tag_id; // @[Decoder.scala 156:31]
  assign valueSelector2_io_reorderBufferValue_valid = io_reorderBuffer_source2_value_valid; // @[Decoder.scala 169:40]
  assign valueSelector2_io_reorderBufferValue_bits = io_reorderBuffer_source2_value_bits; // @[Decoder.scala 169:40]
  assign valueSelector2_io_registerFileValue = io_registerFile_value2; // @[Decoder.scala 170:39]
  assign valueSelector2_io_programCounter = io_instructionFetch_bits_programCounter; // @[Decoder.scala 171:36]
  assign valueSelector2_io_outputCollector_outputs_valid = io_outputCollector_outputs_valid; // @[Decoder.scala 173:37]
  assign valueSelector2_io_outputCollector_outputs_bits_resultType = io_outputCollector_outputs_bits_resultType; // @[Decoder.scala 173:37]
  assign valueSelector2_io_outputCollector_outputs_bits_value = io_outputCollector_outputs_bits_value; // @[Decoder.scala 173:37]
  assign valueSelector2_io_outputCollector_outputs_bits_tag_threadId = io_outputCollector_outputs_bits_tag_threadId; // @[Decoder.scala 173:37]
  assign valueSelector2_io_outputCollector_outputs_bits_tag_id = io_outputCollector_outputs_bits_tag_id; // @[Decoder.scala 173:37]
  assign valueSelector2_io_opcodeFormat = opcodeFormatChecker_io_format; // @[Decoder.scala 172:34]
  assign valueSelector2_io_sourceTag_valid = sourceTagSelector2_io_sourceTag_valid; // @[Decoder.scala 168:31]
  assign valueSelector2_io_sourceTag_tag_threadId = sourceTagSelector2_io_sourceTag_tag_threadId; // @[Decoder.scala 168:31]
  assign valueSelector2_io_sourceTag_tag_id = sourceTagSelector2_io_sourceTag_tag_id; // @[Decoder.scala 168:31]
endmodule
module Decoder_1(
  output        io_instructionFetch_ready,
  input         io_instructionFetch_valid,
  input  [31:0] io_instructionFetch_bits_instruction,
  input  [63:0] io_instructionFetch_bits_programCounter,
  input         io_instructionFetch_bits_wasCompressed,
  output [4:0]  io_reorderBuffer_source1_sourceRegister,
  input         io_reorderBuffer_source1_matchingTag_valid,
  input  [3:0]  io_reorderBuffer_source1_matchingTag_bits_id,
  input         io_reorderBuffer_source1_value_valid,
  input  [63:0] io_reorderBuffer_source1_value_bits,
  output [4:0]  io_reorderBuffer_source2_sourceRegister,
  input         io_reorderBuffer_source2_matchingTag_valid,
  input  [3:0]  io_reorderBuffer_source2_matchingTag_bits_id,
  input         io_reorderBuffer_source2_value_valid,
  input  [63:0] io_reorderBuffer_source2_value_bits,
  output [4:0]  io_reorderBuffer_destination_destinationRegister,
  input  [3:0]  io_reorderBuffer_destination_destinationTag_id,
  output        io_reorderBuffer_destination_storeSign,
  input         io_reorderBuffer_ready,
  output        io_reorderBuffer_valid,
  input         io_outputCollector_outputs_valid,
  input         io_outputCollector_outputs_bits_resultType,
  input  [63:0] io_outputCollector_outputs_bits_value,
  input         io_outputCollector_outputs_bits_tag_threadId,
  input  [3:0]  io_outputCollector_outputs_bits_tag_id,
  output [4:0]  io_registerFile_sourceRegister1,
  output [4:0]  io_registerFile_sourceRegister2,
  input  [63:0] io_registerFile_value1,
  input  [63:0] io_registerFile_value2,
  input         io_reservationStation_ready,
  output [6:0]  io_reservationStation_entry_opcode,
  output [2:0]  io_reservationStation_entry_function3,
  output [11:0] io_reservationStation_entry_immediateOrFunction7,
  output        io_reservationStation_entry_sourceTag1_threadId,
  output [3:0]  io_reservationStation_entry_sourceTag1_id,
  output        io_reservationStation_entry_ready1,
  output [63:0] io_reservationStation_entry_value1,
  output        io_reservationStation_entry_sourceTag2_threadId,
  output [3:0]  io_reservationStation_entry_sourceTag2_id,
  output        io_reservationStation_entry_ready2,
  output [63:0] io_reservationStation_entry_value2,
  output        io_reservationStation_entry_destinationTag_threadId,
  output [3:0]  io_reservationStation_entry_destinationTag_id,
  output        io_reservationStation_entry_wasCompressed,
  output        io_reservationStation_entry_valid,
  input         io_loadStoreQueue_ready,
  output        io_loadStoreQueue_valid,
  output        io_loadStoreQueue_bits_accessInfo_accessType,
  output        io_loadStoreQueue_bits_accessInfo_signed,
  output [1:0]  io_loadStoreQueue_bits_accessInfo_accessWidth,
  output        io_loadStoreQueue_bits_addressAndLoadResultTag_threadId,
  output [3:0]  io_loadStoreQueue_bits_addressAndLoadResultTag_id,
  output [63:0] io_loadStoreQueue_bits_address,
  output        io_loadStoreQueue_bits_addressValid,
  output        io_loadStoreQueue_bits_storeDataTag_threadId,
  output [3:0]  io_loadStoreQueue_bits_storeDataTag_id,
  output [63:0] io_loadStoreQueue_bits_storeData,
  output        io_loadStoreQueue_bits_storeDataValid,
  input         io_csr_ready,
  output        io_csr_valid,
  output        io_csr_bits_sourceTag_threadId,
  output [3:0]  io_csr_bits_sourceTag_id,
  output [3:0]  io_csr_bits_destinationTag_id,
  output [63:0] io_csr_bits_value,
  output        io_csr_bits_ready,
  output [11:0] io_csr_bits_address,
  output [1:0]  io_csr_bits_csrAccessType
);
  wire [6:0] opcodeFormatChecker_io_opcode; // @[Decoder.scala 78:35]
  wire [2:0] opcodeFormatChecker_io_format; // @[Decoder.scala 78:35]
  wire  sourceTagSelector1_io_reorderBufferDestinationTag_valid; // @[Decoder.scala 126:34]
  wire  sourceTagSelector1_io_reorderBufferDestinationTag_bits_threadId; // @[Decoder.scala 126:34]
  wire [3:0] sourceTagSelector1_io_reorderBufferDestinationTag_bits_id; // @[Decoder.scala 126:34]
  wire  sourceTagSelector1_io_sourceTag_valid; // @[Decoder.scala 126:34]
  wire  sourceTagSelector1_io_sourceTag_tag_threadId; // @[Decoder.scala 126:34]
  wire [3:0] sourceTagSelector1_io_sourceTag_tag_id; // @[Decoder.scala 126:34]
  wire  sourceTagSelector2_io_reorderBufferDestinationTag_valid; // @[Decoder.scala 141:34]
  wire  sourceTagSelector2_io_reorderBufferDestinationTag_bits_threadId; // @[Decoder.scala 141:34]
  wire [3:0] sourceTagSelector2_io_reorderBufferDestinationTag_bits_id; // @[Decoder.scala 141:34]
  wire  sourceTagSelector2_io_sourceTag_valid; // @[Decoder.scala 141:34]
  wire  sourceTagSelector2_io_sourceTag_tag_threadId; // @[Decoder.scala 141:34]
  wire [3:0] sourceTagSelector2_io_sourceTag_tag_id; // @[Decoder.scala 141:34]
  wire  valueSelector1_io_reorderBufferValue_valid; // @[Decoder.scala 155:30]
  wire [63:0] valueSelector1_io_reorderBufferValue_bits; // @[Decoder.scala 155:30]
  wire [63:0] valueSelector1_io_registerFileValue; // @[Decoder.scala 155:30]
  wire  valueSelector1_io_outputCollector_outputs_valid; // @[Decoder.scala 155:30]
  wire  valueSelector1_io_outputCollector_outputs_bits_resultType; // @[Decoder.scala 155:30]
  wire [63:0] valueSelector1_io_outputCollector_outputs_bits_value; // @[Decoder.scala 155:30]
  wire  valueSelector1_io_outputCollector_outputs_bits_tag_threadId; // @[Decoder.scala 155:30]
  wire [3:0] valueSelector1_io_outputCollector_outputs_bits_tag_id; // @[Decoder.scala 155:30]
  wire [63:0] valueSelector1_io_immediateValue; // @[Decoder.scala 155:30]
  wire [2:0] valueSelector1_io_opcodeFormat; // @[Decoder.scala 155:30]
  wire  valueSelector1_io_sourceTag_valid; // @[Decoder.scala 155:30]
  wire  valueSelector1_io_sourceTag_tag_threadId; // @[Decoder.scala 155:30]
  wire [3:0] valueSelector1_io_sourceTag_tag_id; // @[Decoder.scala 155:30]
  wire  valueSelector1_io_value_valid; // @[Decoder.scala 155:30]
  wire [63:0] valueSelector1_io_value_bits; // @[Decoder.scala 155:30]
  wire  valueSelector2_io_reorderBufferValue_valid; // @[Decoder.scala 167:30]
  wire [63:0] valueSelector2_io_reorderBufferValue_bits; // @[Decoder.scala 167:30]
  wire [63:0] valueSelector2_io_registerFileValue; // @[Decoder.scala 167:30]
  wire [63:0] valueSelector2_io_programCounter; // @[Decoder.scala 167:30]
  wire  valueSelector2_io_outputCollector_outputs_valid; // @[Decoder.scala 167:30]
  wire  valueSelector2_io_outputCollector_outputs_bits_resultType; // @[Decoder.scala 167:30]
  wire [63:0] valueSelector2_io_outputCollector_outputs_bits_value; // @[Decoder.scala 167:30]
  wire  valueSelector2_io_outputCollector_outputs_bits_tag_threadId; // @[Decoder.scala 167:30]
  wire [3:0] valueSelector2_io_outputCollector_outputs_bits_tag_id; // @[Decoder.scala 167:30]
  wire [2:0] valueSelector2_io_opcodeFormat; // @[Decoder.scala 167:30]
  wire  valueSelector2_io_sourceTag_valid; // @[Decoder.scala 167:30]
  wire  valueSelector2_io_sourceTag_tag_threadId; // @[Decoder.scala 167:30]
  wire [3:0] valueSelector2_io_sourceTag_tag_id; // @[Decoder.scala 167:30]
  wire  valueSelector2_io_value_valid; // @[Decoder.scala 167:30]
  wire [63:0] valueSelector2_io_value_bits; // @[Decoder.scala 167:30]
  wire [4:0] instRd = io_instructionFetch_bits_instruction[11:7]; // @[Decoder.scala 46:52]
  wire [4:0] instRs1 = io_instructionFetch_bits_instruction[19:15]; // @[Decoder.scala 47:53]
  wire [4:0] instRs2 = io_instructionFetch_bits_instruction[24:20]; // @[Decoder.scala 48:53]
  wire [2:0] instFunct3 = io_instructionFetch_bits_instruction[14:12]; // @[Decoder.scala 49:56]
  wire [6:0] instFunct7 = io_instructionFetch_bits_instruction[31:25]; // @[Decoder.scala 50:56]
  wire [6:0] instOp = io_instructionFetch_bits_instruction[6:0]; // @[Decoder.scala 51:52]
  wire [11:0] instImmS = {instFunct7,instRd}; // @[Cat.scala 33:92]
  wire [11:0] instImmB = {io_instructionFetch_bits_instruction[31],io_instructionFetch_bits_instruction[7],
    io_instructionFetch_bits_instruction[30:25],io_instructionFetch_bits_instruction[11:8]}; // @[Cat.scala 33:92]
  wire [19:0] instImmU = io_instructionFetch_bits_instruction[31:12]; // @[Decoder.scala 63:54]
  wire [11:0] immIExtended = io_instructionFetch_bits_instruction[31:20]; // @[Decoder.scala 73:14]
  wire [31:0] immUExtended = {instImmU,12'h0}; // @[Decoder.scala 74:47]
  wire [20:0] immJExtended = {io_instructionFetch_bits_instruction[31],io_instructionFetch_bits_instruction[19:12],
    io_instructionFetch_bits_instruction[20],io_instructionFetch_bits_instruction[30:21],1'h0}; // @[Decoder.scala 75:46]
  wire  _destinationIsValid_T = opcodeFormatChecker_io_format == 3'h0; // @[Decoder.scala 82:58]
  wire  _destinationIsValid_T_1 = opcodeFormatChecker_io_format == 3'h1; // @[Decoder.scala 83:35]
  wire  _destinationIsValid_T_2 = opcodeFormatChecker_io_format == 3'h0 | _destinationIsValid_T_1; // @[Decoder.scala 82:64]
  wire  _destinationIsValid_T_3 = opcodeFormatChecker_io_format == 3'h4; // @[Decoder.scala 84:35]
  wire  _destinationIsValid_T_4 = _destinationIsValid_T_2 | _destinationIsValid_T_3; // @[Decoder.scala 83:41]
  wire  _destinationIsValid_T_5 = opcodeFormatChecker_io_format == 3'h2; // @[Decoder.scala 85:35]
  wire  destinationIsValid = _destinationIsValid_T_4 | _destinationIsValid_T_5; // @[Decoder.scala 84:41]
  wire  _source1IsValid_T_3 = opcodeFormatChecker_io_format == 3'h3; // @[Decoder.scala 90:35]
  wire  _source1IsValid_T_4 = _destinationIsValid_T_2 | _source1IsValid_T_3; // @[Decoder.scala 89:41]
  wire  _source1IsValid_T_5 = opcodeFormatChecker_io_format == 3'h5; // @[Decoder.scala 91:35]
  wire  source1IsValid = _source1IsValid_T_4 | _source1IsValid_T_5; // @[Decoder.scala 90:41]
  wire  _source2IsValid_T_2 = _destinationIsValid_T | _source1IsValid_T_3; // @[Decoder.scala 94:60]
  wire  source2IsValid = _source2IsValid_T_2 | _source1IsValid_T_5; // @[Decoder.scala 95:41]
  wire  _io_reorderBuffer_destination_storeSign_T = instOp == 7'h23; // @[Decoder.scala 106:52]
  wire [2:0] _valueSelector1_io_immediateValue_T = opcodeFormatChecker_io_format; // @[Decoder.scala 162:35]
  wire [31:0] _valueSelector1_io_immediateValue_T_4 = 3'h4 == _valueSelector1_io_immediateValue_T ? $signed(immUExtended
    ) : $signed(32'sh0); // @[Mux.scala 81:58]
  wire [31:0] _valueSelector1_io_immediateValue_T_6 = 3'h2 == _valueSelector1_io_immediateValue_T ? $signed({{11{
    immJExtended[20]}},immJExtended}) : $signed(_valueSelector1_io_immediateValue_T_4); // @[Mux.scala 81:58]
  wire  _io_reorderBuffer_valid_T = io_instructionFetch_ready & io_instructionFetch_valid; // @[Decoder.scala 194:55]
  wire [6:0] _io_reservationStation_entry_valid_T_1 = instOp & 7'h5f; // @[Decoder.scala 197:14]
  wire  _io_reservationStation_entry_valid_T_2 = 7'h3 == _io_reservationStation_entry_valid_T_1; // @[Decoder.scala 197:14]
  wire  _io_reservationStation_entry_valid_T_3 = _io_reservationStation_entry_valid_T_2 & valueSelector1_io_value_valid; // @[Decoder.scala 199:7]
  wire  _io_reservationStation_entry_valid_T_4 = ~_io_reservationStation_entry_valid_T_3; // @[Decoder.scala 197:5]
  wire  _io_reservationStation_entry_valid_T_5 = _io_reorderBuffer_valid_T & _io_reservationStation_entry_valid_T_4; // @[Decoder.scala 196:31]
  wire [11:0] _io_reservationStation_entry_immediateOrFunction7_T_2 = {instFunct7,5'h0}; // @[Cat.scala 33:92]
  wire [11:0] _io_reservationStation_entry_immediateOrFunction7_T_6 = io_instructionFetch_bits_instruction[31:20]; // @[Decoder.scala 212:32]
  wire [11:0] _io_reservationStation_entry_immediateOrFunction7_T_8 = 3'h0 == _valueSelector1_io_immediateValue_T ?
    _io_reservationStation_entry_immediateOrFunction7_T_2 : 12'h0; // @[Mux.scala 81:58]
  wire [11:0] _io_reservationStation_entry_immediateOrFunction7_T_10 = 3'h3 == _valueSelector1_io_immediateValue_T ?
    instImmS : _io_reservationStation_entry_immediateOrFunction7_T_8; // @[Mux.scala 81:58]
  wire [11:0] _io_reservationStation_entry_immediateOrFunction7_T_12 = 3'h5 == _valueSelector1_io_immediateValue_T ?
    instImmB : _io_reservationStation_entry_immediateOrFunction7_T_10; // @[Mux.scala 81:58]
  wire  _io_loadStoreQueue_valid_T_2 = io_loadStoreQueue_ready & _io_reservationStation_entry_valid_T_2; // @[Decoder.scala 233:54]
  wire  _io_loadStoreQueue_bits_accessInfo_w_accessWidth_T_3 = instFunct3[1:0] == 2'h1; // @[MemoryAccessWidth.scala 13:23]
  wire  _io_loadStoreQueue_bits_accessInfo_w_accessWidth_T_5 = instFunct3[1:0] == 2'h2; // @[MemoryAccessWidth.scala 14:23]
  wire  _io_loadStoreQueue_bits_accessInfo_w_accessWidth_T_7 = instFunct3[1:0] == 2'h3; // @[MemoryAccessWidth.scala 15:23]
  wire [1:0] _io_loadStoreQueue_bits_accessInfo_w_accessWidth_T_13 =
    _io_loadStoreQueue_bits_accessInfo_w_accessWidth_T_5 ? 2'h2 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_loadStoreQueue_bits_accessInfo_w_accessWidth_T_15 =
    _io_loadStoreQueue_bits_accessInfo_w_accessWidth_T_7 ? 2'h3 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _GEN_27 = {{1'd0}, _io_loadStoreQueue_bits_accessInfo_w_accessWidth_T_3}; // @[Mux.scala 27:73]
  wire [1:0] _io_loadStoreQueue_bits_accessInfo_w_accessWidth_T_17 = _GEN_27 |
    _io_loadStoreQueue_bits_accessInfo_w_accessWidth_T_13; // @[Mux.scala 27:73]
  wire [11:0] _io_loadStoreQueue_bits_address_T_2 = {instFunct7,instRd}; // @[Decoder.scala 245:16]
  wire [11:0] _io_loadStoreQueue_bits_address_T_4 = _io_reorderBuffer_destination_storeSign_T ? $signed(
    _io_loadStoreQueue_bits_address_T_2) : $signed(immIExtended); // @[Decoder.scala 243:81]
  wire [63:0] _GEN_28 = {{52{_io_loadStoreQueue_bits_address_T_4[11]}},_io_loadStoreQueue_bits_address_T_4}; // @[Decoder.scala 243:76]
  OpcodeFormatChecker opcodeFormatChecker ( // @[Decoder.scala 78:35]
    .io_opcode(opcodeFormatChecker_io_opcode),
    .io_format(opcodeFormatChecker_io_format)
  );
  SourceTagSelector sourceTagSelector1 ( // @[Decoder.scala 126:34]
    .io_reorderBufferDestinationTag_valid(sourceTagSelector1_io_reorderBufferDestinationTag_valid),
    .io_reorderBufferDestinationTag_bits_threadId(sourceTagSelector1_io_reorderBufferDestinationTag_bits_threadId),
    .io_reorderBufferDestinationTag_bits_id(sourceTagSelector1_io_reorderBufferDestinationTag_bits_id),
    .io_sourceTag_valid(sourceTagSelector1_io_sourceTag_valid),
    .io_sourceTag_tag_threadId(sourceTagSelector1_io_sourceTag_tag_threadId),
    .io_sourceTag_tag_id(sourceTagSelector1_io_sourceTag_tag_id)
  );
  SourceTagSelector sourceTagSelector2 ( // @[Decoder.scala 141:34]
    .io_reorderBufferDestinationTag_valid(sourceTagSelector2_io_reorderBufferDestinationTag_valid),
    .io_reorderBufferDestinationTag_bits_threadId(sourceTagSelector2_io_reorderBufferDestinationTag_bits_threadId),
    .io_reorderBufferDestinationTag_bits_id(sourceTagSelector2_io_reorderBufferDestinationTag_bits_id),
    .io_sourceTag_valid(sourceTagSelector2_io_sourceTag_valid),
    .io_sourceTag_tag_threadId(sourceTagSelector2_io_sourceTag_tag_threadId),
    .io_sourceTag_tag_id(sourceTagSelector2_io_sourceTag_tag_id)
  );
  ValueSelector1 valueSelector1 ( // @[Decoder.scala 155:30]
    .io_reorderBufferValue_valid(valueSelector1_io_reorderBufferValue_valid),
    .io_reorderBufferValue_bits(valueSelector1_io_reorderBufferValue_bits),
    .io_registerFileValue(valueSelector1_io_registerFileValue),
    .io_outputCollector_outputs_valid(valueSelector1_io_outputCollector_outputs_valid),
    .io_outputCollector_outputs_bits_resultType(valueSelector1_io_outputCollector_outputs_bits_resultType),
    .io_outputCollector_outputs_bits_value(valueSelector1_io_outputCollector_outputs_bits_value),
    .io_outputCollector_outputs_bits_tag_threadId(valueSelector1_io_outputCollector_outputs_bits_tag_threadId),
    .io_outputCollector_outputs_bits_tag_id(valueSelector1_io_outputCollector_outputs_bits_tag_id),
    .io_immediateValue(valueSelector1_io_immediateValue),
    .io_opcodeFormat(valueSelector1_io_opcodeFormat),
    .io_sourceTag_valid(valueSelector1_io_sourceTag_valid),
    .io_sourceTag_tag_threadId(valueSelector1_io_sourceTag_tag_threadId),
    .io_sourceTag_tag_id(valueSelector1_io_sourceTag_tag_id),
    .io_value_valid(valueSelector1_io_value_valid),
    .io_value_bits(valueSelector1_io_value_bits)
  );
  ValueSelector2 valueSelector2 ( // @[Decoder.scala 167:30]
    .io_reorderBufferValue_valid(valueSelector2_io_reorderBufferValue_valid),
    .io_reorderBufferValue_bits(valueSelector2_io_reorderBufferValue_bits),
    .io_registerFileValue(valueSelector2_io_registerFileValue),
    .io_programCounter(valueSelector2_io_programCounter),
    .io_outputCollector_outputs_valid(valueSelector2_io_outputCollector_outputs_valid),
    .io_outputCollector_outputs_bits_resultType(valueSelector2_io_outputCollector_outputs_bits_resultType),
    .io_outputCollector_outputs_bits_value(valueSelector2_io_outputCollector_outputs_bits_value),
    .io_outputCollector_outputs_bits_tag_threadId(valueSelector2_io_outputCollector_outputs_bits_tag_threadId),
    .io_outputCollector_outputs_bits_tag_id(valueSelector2_io_outputCollector_outputs_bits_tag_id),
    .io_opcodeFormat(valueSelector2_io_opcodeFormat),
    .io_sourceTag_valid(valueSelector2_io_sourceTag_valid),
    .io_sourceTag_tag_threadId(valueSelector2_io_sourceTag_tag_threadId),
    .io_sourceTag_tag_id(valueSelector2_io_sourceTag_tag_id),
    .io_value_valid(valueSelector2_io_value_valid),
    .io_value_bits(valueSelector2_io_value_bits)
  );
  assign io_instructionFetch_ready = io_reservationStation_ready & io_reorderBuffer_ready & io_loadStoreQueue_ready &
    io_csr_ready; // @[Decoder.scala 192:113]
  assign io_reorderBuffer_source1_sourceRegister = source1IsValid ? instRs1 : 5'h0; // @[Decoder.scala 99:49]
  assign io_reorderBuffer_source2_sourceRegister = source2IsValid ? instRs2 : 5'h0; // @[Decoder.scala 100:49]
  assign io_reorderBuffer_destination_destinationRegister = destinationIsValid ? instRd : 5'h0; // @[Decoder.scala 101:58]
  assign io_reorderBuffer_destination_storeSign = instOp == 7'h23; // @[Decoder.scala 106:52]
  assign io_reorderBuffer_valid = io_instructionFetch_ready & io_instructionFetch_valid; // @[Decoder.scala 194:55]
  assign io_registerFile_sourceRegister1 = io_instructionFetch_bits_instruction[19:15]; // @[Decoder.scala 47:53]
  assign io_registerFile_sourceRegister2 = io_instructionFetch_bits_instruction[24:20]; // @[Decoder.scala 48:53]
  assign io_reservationStation_entry_opcode = io_instructionFetch_bits_instruction[6:0]; // @[Decoder.scala 51:52]
  assign io_reservationStation_entry_function3 = io_instructionFetch_bits_instruction[14:12]; // @[Decoder.scala 49:56]
  assign io_reservationStation_entry_immediateOrFunction7 = 3'h1 == _valueSelector1_io_immediateValue_T ?
    _io_reservationStation_entry_immediateOrFunction7_T_6 : _io_reservationStation_entry_immediateOrFunction7_T_12; // @[Mux.scala 81:58]
  assign io_reservationStation_entry_sourceTag1_threadId = valueSelector1_io_value_valid |
    sourceTagSelector1_io_sourceTag_tag_threadId; // @[Decoder.scala 216:23]
  assign io_reservationStation_entry_sourceTag1_id = valueSelector1_io_value_valid ? 4'h0 :
    sourceTagSelector1_io_sourceTag_tag_id; // @[Decoder.scala 216:23]
  assign io_reservationStation_entry_ready1 = valueSelector1_io_value_valid; // @[Decoder.scala 226:13]
  assign io_reservationStation_entry_value1 = valueSelector1_io_value_bits; // @[Decoder.scala 228:13]
  assign io_reservationStation_entry_sourceTag2_threadId = valueSelector2_io_value_valid |
    sourceTagSelector2_io_sourceTag_tag_threadId; // @[Decoder.scala 221:23]
  assign io_reservationStation_entry_sourceTag2_id = valueSelector2_io_value_valid ? 4'h0 :
    sourceTagSelector2_io_sourceTag_tag_id; // @[Decoder.scala 221:23]
  assign io_reservationStation_entry_ready2 = valueSelector2_io_value_valid; // @[Decoder.scala 227:13]
  assign io_reservationStation_entry_value2 = valueSelector2_io_value_bits; // @[Decoder.scala 229:13]
  assign io_reservationStation_entry_destinationTag_threadId = 1'h1; // @[Decoder.scala 215:21]
  assign io_reservationStation_entry_destinationTag_id = io_reorderBuffer_destination_destinationTag_id; // @[Decoder.scala 215:21]
  assign io_reservationStation_entry_wasCompressed = io_instructionFetch_bits_wasCompressed; // @[Decoder.scala 230:20]
  assign io_reservationStation_entry_valid = _io_reservationStation_entry_valid_T_5 & instOp != 7'h73; // @[Decoder.scala 199:41]
  assign io_loadStoreQueue_valid = _io_loadStoreQueue_valid_T_2 & io_instructionFetch_ready & io_instructionFetch_valid; // @[Decoder.scala 235:34]
  assign io_loadStoreQueue_bits_accessInfo_accessType = ~instOp[5]; // @[MemoryAccessType.scala 15:20]
  assign io_loadStoreQueue_bits_accessInfo_signed = ~instFunct3[2]; // @[MemoryAccessInfo.scala 15:17]
  assign io_loadStoreQueue_bits_accessInfo_accessWidth = _io_loadStoreQueue_bits_accessInfo_w_accessWidth_T_17 |
    _io_loadStoreQueue_bits_accessInfo_w_accessWidth_T_15; // @[Mux.scala 27:73]
  assign io_loadStoreQueue_bits_addressAndLoadResultTag_threadId = io_reservationStation_entry_destinationTag_threadId; // @[Decoder.scala 239:33 241:52]
  assign io_loadStoreQueue_bits_addressAndLoadResultTag_id = io_reservationStation_entry_destinationTag_id; // @[Decoder.scala 239:33 241:52]
  assign io_loadStoreQueue_bits_address = $signed(valueSelector1_io_value_bits) + $signed(_GEN_28); // @[Decoder.scala 247:8]
  assign io_loadStoreQueue_bits_addressValid = valueSelector1_io_value_valid; // @[Decoder.scala 239:33 242:41]
  assign io_loadStoreQueue_bits_storeDataTag_threadId = _io_reorderBuffer_destination_storeSign_T ?
    valueSelector2_io_sourceTag_tag_threadId : 1'h1; // @[Decoder.scala 248:28 249:43 253:43]
  assign io_loadStoreQueue_bits_storeDataTag_id = _io_reorderBuffer_destination_storeSign_T ?
    valueSelector2_io_sourceTag_tag_id : 4'h0; // @[Decoder.scala 248:28 249:43 253:43]
  assign io_loadStoreQueue_bits_storeData = _io_reorderBuffer_destination_storeSign_T ? valueSelector2_io_value_bits : 64'h0
    ; // @[Decoder.scala 248:28 250:40 254:40]
  assign io_loadStoreQueue_bits_storeDataValid = _io_reorderBuffer_destination_storeSign_T ?
    valueSelector2_io_value_valid : 1'h1; // @[Decoder.scala 248:28 251:45 255:45]
  assign io_csr_valid = io_csr_ready & io_instructionFetch_ready & io_instructionFetch_valid & 7'h73 == instOp &
    instFunct3 != 3'h0; // @[Decoder.scala 261:117]
  assign io_csr_bits_sourceTag_threadId = valueSelector1_io_sourceTag_tag_threadId; // @[Decoder.scala 263:22 274:27]
  assign io_csr_bits_sourceTag_id = valueSelector1_io_sourceTag_tag_id; // @[Decoder.scala 263:22 274:27]
  assign io_csr_bits_destinationTag_id = io_reorderBuffer_destination_destinationTag_id; // @[Decoder.scala 263:22 285:32]
  assign io_csr_bits_value = instFunct3[2] ? {{59'd0}, instRs1} : valueSelector1_io_value_bits; // @[Decoder.scala 275:29]
  assign io_csr_bits_ready = instFunct3[2] | valueSelector1_io_value_valid; // @[Decoder.scala 280:29]
  assign io_csr_bits_address = io_instructionFetch_bits_instruction[31:20]; // @[Decoder.scala 52:54]
  assign io_csr_bits_csrAccessType = 2'h3 == instFunct3[1:0] ? 2'h2 : {{1'd0}, 2'h2 == instFunct3[1:0]}; // @[Mux.scala 81:58]
  assign opcodeFormatChecker_io_opcode = io_instructionFetch_bits_instruction[6:0]; // @[Decoder.scala 51:52]
  assign sourceTagSelector1_io_reorderBufferDestinationTag_valid = io_reorderBuffer_source1_matchingTag_valid; // @[Decoder.scala 127:53]
  assign sourceTagSelector1_io_reorderBufferDestinationTag_bits_threadId = 1'h1; // @[Decoder.scala 127:53]
  assign sourceTagSelector1_io_reorderBufferDestinationTag_bits_id = io_reorderBuffer_source1_matchingTag_bits_id; // @[Decoder.scala 127:53]
  assign sourceTagSelector2_io_reorderBufferDestinationTag_valid = io_reorderBuffer_source2_matchingTag_valid; // @[Decoder.scala 142:53]
  assign sourceTagSelector2_io_reorderBufferDestinationTag_bits_threadId = 1'h1; // @[Decoder.scala 142:53]
  assign sourceTagSelector2_io_reorderBufferDestinationTag_bits_id = io_reorderBuffer_source2_matchingTag_bits_id; // @[Decoder.scala 142:53]
  assign valueSelector1_io_reorderBufferValue_valid = io_reorderBuffer_source1_value_valid; // @[Decoder.scala 157:40]
  assign valueSelector1_io_reorderBufferValue_bits = io_reorderBuffer_source1_value_bits; // @[Decoder.scala 157:40]
  assign valueSelector1_io_registerFileValue = io_registerFile_value1; // @[Decoder.scala 158:39]
  assign valueSelector1_io_outputCollector_outputs_valid = io_outputCollector_outputs_valid; // @[Decoder.scala 159:37]
  assign valueSelector1_io_outputCollector_outputs_bits_resultType = io_outputCollector_outputs_bits_resultType; // @[Decoder.scala 159:37]
  assign valueSelector1_io_outputCollector_outputs_bits_value = io_outputCollector_outputs_bits_value; // @[Decoder.scala 159:37]
  assign valueSelector1_io_outputCollector_outputs_bits_tag_threadId = io_outputCollector_outputs_bits_tag_threadId; // @[Decoder.scala 159:37]
  assign valueSelector1_io_outputCollector_outputs_bits_tag_id = io_outputCollector_outputs_bits_tag_id; // @[Decoder.scala 159:37]
  assign valueSelector1_io_immediateValue = {{32{_valueSelector1_io_immediateValue_T_6[31]}},
    _valueSelector1_io_immediateValue_T_6}; // @[Decoder.scala 161:36]
  assign valueSelector1_io_opcodeFormat = opcodeFormatChecker_io_format; // @[Decoder.scala 160:34]
  assign valueSelector1_io_sourceTag_valid = sourceTagSelector1_io_sourceTag_valid; // @[Decoder.scala 156:31]
  assign valueSelector1_io_sourceTag_tag_threadId = sourceTagSelector1_io_sourceTag_tag_threadId; // @[Decoder.scala 156:31]
  assign valueSelector1_io_sourceTag_tag_id = sourceTagSelector1_io_sourceTag_tag_id; // @[Decoder.scala 156:31]
  assign valueSelector2_io_reorderBufferValue_valid = io_reorderBuffer_source2_value_valid; // @[Decoder.scala 169:40]
  assign valueSelector2_io_reorderBufferValue_bits = io_reorderBuffer_source2_value_bits; // @[Decoder.scala 169:40]
  assign valueSelector2_io_registerFileValue = io_registerFile_value2; // @[Decoder.scala 170:39]
  assign valueSelector2_io_programCounter = io_instructionFetch_bits_programCounter; // @[Decoder.scala 171:36]
  assign valueSelector2_io_outputCollector_outputs_valid = io_outputCollector_outputs_valid; // @[Decoder.scala 173:37]
  assign valueSelector2_io_outputCollector_outputs_bits_resultType = io_outputCollector_outputs_bits_resultType; // @[Decoder.scala 173:37]
  assign valueSelector2_io_outputCollector_outputs_bits_value = io_outputCollector_outputs_bits_value; // @[Decoder.scala 173:37]
  assign valueSelector2_io_outputCollector_outputs_bits_tag_threadId = io_outputCollector_outputs_bits_tag_threadId; // @[Decoder.scala 173:37]
  assign valueSelector2_io_outputCollector_outputs_bits_tag_id = io_outputCollector_outputs_bits_tag_id; // @[Decoder.scala 173:37]
  assign valueSelector2_io_opcodeFormat = opcodeFormatChecker_io_format; // @[Decoder.scala 172:34]
  assign valueSelector2_io_sourceTag_valid = sourceTagSelector2_io_sourceTag_valid; // @[Decoder.scala 168:31]
  assign valueSelector2_io_sourceTag_tag_threadId = sourceTagSelector2_io_sourceTag_tag_threadId; // @[Decoder.scala 168:31]
  assign valueSelector2_io_sourceTag_tag_id = sourceTagSelector2_io_sourceTag_tag_id; // @[Decoder.scala 168:31]
endmodule
module B4RRArbiter_1(
  input         clock,
  input         reset,
  output        io_in_0_ready,
  input         io_in_0_valid,
  input         io_in_0_bits_destinationTag_threadId,
  input  [3:0]  io_in_0_bits_destinationTag_id,
  input  [63:0] io_in_0_bits_value1,
  input  [63:0] io_in_0_bits_value2,
  input  [2:0]  io_in_0_bits_function3,
  input  [11:0] io_in_0_bits_immediateOrFunction7,
  input  [6:0]  io_in_0_bits_opcode,
  input         io_in_0_bits_wasCompressed,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input         io_in_1_bits_destinationTag_threadId,
  input  [3:0]  io_in_1_bits_destinationTag_id,
  input  [63:0] io_in_1_bits_value1,
  input  [63:0] io_in_1_bits_value2,
  input  [2:0]  io_in_1_bits_function3,
  input  [11:0] io_in_1_bits_immediateOrFunction7,
  input  [6:0]  io_in_1_bits_opcode,
  input         io_in_1_bits_wasCompressed,
  output        io_in_2_ready,
  input         io_in_2_valid,
  input         io_in_2_bits_destinationTag_threadId,
  input  [3:0]  io_in_2_bits_destinationTag_id,
  input  [63:0] io_in_2_bits_value1,
  input  [63:0] io_in_2_bits_value2,
  input  [2:0]  io_in_2_bits_function3,
  input  [11:0] io_in_2_bits_immediateOrFunction7,
  input  [6:0]  io_in_2_bits_opcode,
  input         io_in_2_bits_wasCompressed,
  output        io_in_3_ready,
  input         io_in_3_valid,
  input         io_in_3_bits_destinationTag_threadId,
  input  [3:0]  io_in_3_bits_destinationTag_id,
  input  [63:0] io_in_3_bits_value1,
  input  [63:0] io_in_3_bits_value2,
  input  [2:0]  io_in_3_bits_function3,
  input  [11:0] io_in_3_bits_immediateOrFunction7,
  input  [6:0]  io_in_3_bits_opcode,
  input         io_in_3_bits_wasCompressed,
  input         io_out_ready,
  output        io_out_valid,
  output        io_out_bits_destinationTag_threadId,
  output [3:0]  io_out_bits_destinationTag_id,
  output [63:0] io_out_bits_value1,
  output [63:0] io_out_bits_value2,
  output [2:0]  io_out_bits_function3,
  output [11:0] io_out_bits_immediateOrFunction7,
  output [6:0]  io_out_bits_opcode,
  output        io_out_bits_wasCompressed,
  output [1:0]  io_chosen
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  _GEN_1 = 2'h1 == io_chosen ? io_in_1_valid : io_in_0_valid; // @[Arbitar.scala 59:{16,16}]
  wire  _GEN_2 = 2'h2 == io_chosen ? io_in_2_valid : _GEN_1; // @[Arbitar.scala 59:{16,16}]
  wire  _GEN_5 = 2'h1 == io_chosen ? io_in_1_bits_destinationTag_threadId : io_in_0_bits_destinationTag_threadId; // @[Arbitar.scala 60:{15,15}]
  wire  _GEN_6 = 2'h2 == io_chosen ? io_in_2_bits_destinationTag_threadId : _GEN_5; // @[Arbitar.scala 60:{15,15}]
  wire [3:0] _GEN_9 = 2'h1 == io_chosen ? io_in_1_bits_destinationTag_id : io_in_0_bits_destinationTag_id; // @[Arbitar.scala 60:{15,15}]
  wire [3:0] _GEN_10 = 2'h2 == io_chosen ? io_in_2_bits_destinationTag_id : _GEN_9; // @[Arbitar.scala 60:{15,15}]
  wire [63:0] _GEN_13 = 2'h1 == io_chosen ? io_in_1_bits_value1 : io_in_0_bits_value1; // @[Arbitar.scala 60:{15,15}]
  wire [63:0] _GEN_14 = 2'h2 == io_chosen ? io_in_2_bits_value1 : _GEN_13; // @[Arbitar.scala 60:{15,15}]
  wire [63:0] _GEN_17 = 2'h1 == io_chosen ? io_in_1_bits_value2 : io_in_0_bits_value2; // @[Arbitar.scala 60:{15,15}]
  wire [63:0] _GEN_18 = 2'h2 == io_chosen ? io_in_2_bits_value2 : _GEN_17; // @[Arbitar.scala 60:{15,15}]
  wire [2:0] _GEN_21 = 2'h1 == io_chosen ? io_in_1_bits_function3 : io_in_0_bits_function3; // @[Arbitar.scala 60:{15,15}]
  wire [2:0] _GEN_22 = 2'h2 == io_chosen ? io_in_2_bits_function3 : _GEN_21; // @[Arbitar.scala 60:{15,15}]
  wire [11:0] _GEN_25 = 2'h1 == io_chosen ? io_in_1_bits_immediateOrFunction7 : io_in_0_bits_immediateOrFunction7; // @[Arbitar.scala 60:{15,15}]
  wire [11:0] _GEN_26 = 2'h2 == io_chosen ? io_in_2_bits_immediateOrFunction7 : _GEN_25; // @[Arbitar.scala 60:{15,15}]
  wire [6:0] _GEN_29 = 2'h1 == io_chosen ? io_in_1_bits_opcode : io_in_0_bits_opcode; // @[Arbitar.scala 60:{15,15}]
  wire [6:0] _GEN_30 = 2'h2 == io_chosen ? io_in_2_bits_opcode : _GEN_29; // @[Arbitar.scala 60:{15,15}]
  wire  _GEN_33 = 2'h1 == io_chosen ? io_in_1_bits_wasCompressed : io_in_0_bits_wasCompressed; // @[Arbitar.scala 60:{15,15}]
  wire  _GEN_34 = 2'h2 == io_chosen ? io_in_2_bits_wasCompressed : _GEN_33; // @[Arbitar.scala 60:{15,15}]
  wire  _ctrl_validMask_grantMask_lastGrant_T = io_out_ready & io_out_valid; // @[Decoupled.scala 51:35]
  reg [1:0] lastGrant; // @[Reg.scala 35:20]
  wire  grantMask_1 = 2'h1 > lastGrant; // @[Arbitar.scala 89:49]
  wire  grantMask_2 = 2'h2 > lastGrant; // @[Arbitar.scala 89:49]
  wire  grantMask_3 = 2'h3 > lastGrant; // @[Arbitar.scala 89:49]
  wire  validMask_1 = io_in_1_valid & grantMask_1; // @[Arbitar.scala 91:57]
  wire  validMask_2 = io_in_2_valid & grantMask_2; // @[Arbitar.scala 91:57]
  wire  validMask_3 = io_in_3_valid & grantMask_3; // @[Arbitar.scala 91:57]
  wire  ctrl_2 = ~validMask_1; // @[Arbitar.scala 44:78]
  wire  ctrl_3 = ~(validMask_1 | validMask_2); // @[Arbitar.scala 44:78]
  wire  ctrl_4 = ~(validMask_1 | validMask_2 | validMask_3); // @[Arbitar.scala 44:78]
  wire  ctrl_5 = ~(validMask_1 | validMask_2 | validMask_3 | io_in_0_valid); // @[Arbitar.scala 44:78]
  wire  ctrl_6 = ~(validMask_1 | validMask_2 | validMask_3 | io_in_0_valid | io_in_1_valid); // @[Arbitar.scala 44:78]
  wire  ctrl_7 = ~(validMask_1 | validMask_2 | validMask_3 | io_in_0_valid | io_in_1_valid | io_in_2_valid); // @[Arbitar.scala 44:78]
  wire  _T_3 = grantMask_1 | ctrl_5; // @[Arbitar.scala 97:50]
  wire  _T_5 = ctrl_2 & grantMask_2 | ctrl_6; // @[Arbitar.scala 97:50]
  wire  _T_7 = ctrl_3 & grantMask_3 | ctrl_7; // @[Arbitar.scala 97:50]
  wire [1:0] _GEN_37 = io_in_2_valid ? 2'h2 : 2'h3; // @[Arbitar.scala 102:{26,35} 100:41]
  wire [1:0] _GEN_38 = io_in_1_valid ? 2'h1 : _GEN_37; // @[Arbitar.scala 102:{26,35}]
  wire [1:0] _GEN_39 = io_in_0_valid ? 2'h0 : _GEN_38; // @[Arbitar.scala 102:{26,35}]
  wire [1:0] _GEN_40 = validMask_3 ? 2'h3 : _GEN_39; // @[Arbitar.scala 104:{24,33}]
  wire [1:0] _GEN_41 = validMask_2 ? 2'h2 : _GEN_40; // @[Arbitar.scala 104:{24,33}]
  assign io_in_0_ready = ctrl_4 & io_out_ready; // @[Arbitar.scala 78:21]
  assign io_in_1_ready = _T_3 & io_out_ready; // @[Arbitar.scala 78:21]
  assign io_in_2_ready = _T_5 & io_out_ready; // @[Arbitar.scala 78:21]
  assign io_in_3_ready = _T_7 & io_out_ready; // @[Arbitar.scala 78:21]
  assign io_out_valid = 2'h3 == io_chosen ? io_in_3_valid : _GEN_2; // @[Arbitar.scala 59:{16,16}]
  assign io_out_bits_destinationTag_threadId = 2'h3 == io_chosen ? io_in_3_bits_destinationTag_threadId : _GEN_6; // @[Arbitar.scala 60:{15,15}]
  assign io_out_bits_destinationTag_id = 2'h3 == io_chosen ? io_in_3_bits_destinationTag_id : _GEN_10; // @[Arbitar.scala 60:{15,15}]
  assign io_out_bits_value1 = 2'h3 == io_chosen ? io_in_3_bits_value1 : _GEN_14; // @[Arbitar.scala 60:{15,15}]
  assign io_out_bits_value2 = 2'h3 == io_chosen ? io_in_3_bits_value2 : _GEN_18; // @[Arbitar.scala 60:{15,15}]
  assign io_out_bits_function3 = 2'h3 == io_chosen ? io_in_3_bits_function3 : _GEN_22; // @[Arbitar.scala 60:{15,15}]
  assign io_out_bits_immediateOrFunction7 = 2'h3 == io_chosen ? io_in_3_bits_immediateOrFunction7 : _GEN_26; // @[Arbitar.scala 60:{15,15}]
  assign io_out_bits_opcode = 2'h3 == io_chosen ? io_in_3_bits_opcode : _GEN_30; // @[Arbitar.scala 60:{15,15}]
  assign io_out_bits_wasCompressed = 2'h3 == io_chosen ? io_in_3_bits_wasCompressed : _GEN_34; // @[Arbitar.scala 60:{15,15}]
  assign io_chosen = validMask_1 ? 2'h1 : _GEN_41; // @[Arbitar.scala 104:{24,33}]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 35:20]
      lastGrant <= 2'h0; // @[Reg.scala 35:20]
    end else if (_ctrl_validMask_grantMask_lastGrant_T) begin // @[Reg.scala 36:18]
      lastGrant <= io_chosen; // @[Reg.scala 36:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  lastGrant = _RAND_0[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ReservationStation(
  input         clock,
  input         reset,
  input         io_collectedOutput_0_outputs_valid,
  input         io_collectedOutput_0_outputs_bits_resultType,
  input  [63:0] io_collectedOutput_0_outputs_bits_value,
  input         io_collectedOutput_0_outputs_bits_tag_threadId,
  input  [3:0]  io_collectedOutput_0_outputs_bits_tag_id,
  input         io_collectedOutput_1_outputs_valid,
  input         io_collectedOutput_1_outputs_bits_resultType,
  input  [63:0] io_collectedOutput_1_outputs_bits_value,
  input         io_collectedOutput_1_outputs_bits_tag_threadId,
  input  [3:0]  io_collectedOutput_1_outputs_bits_tag_id,
  input         io_executor_0_ready,
  output        io_executor_0_valid,
  output        io_executor_0_bits_destinationTag_threadId,
  output [3:0]  io_executor_0_bits_destinationTag_id,
  output [63:0] io_executor_0_bits_value1,
  output [63:0] io_executor_0_bits_value2,
  output [2:0]  io_executor_0_bits_function3,
  output [11:0] io_executor_0_bits_immediateOrFunction7,
  output [6:0]  io_executor_0_bits_opcode,
  output        io_executor_0_bits_wasCompressed,
  input         io_executor_1_ready,
  output        io_executor_1_valid,
  output        io_executor_1_bits_destinationTag_threadId,
  output [3:0]  io_executor_1_bits_destinationTag_id,
  output [63:0] io_executor_1_bits_value1,
  output [63:0] io_executor_1_bits_value2,
  output [2:0]  io_executor_1_bits_function3,
  output [11:0] io_executor_1_bits_immediateOrFunction7,
  output [6:0]  io_executor_1_bits_opcode,
  output        io_executor_1_bits_wasCompressed,
  output        io_decoder_0_ready,
  input  [6:0]  io_decoder_0_entry_opcode,
  input  [2:0]  io_decoder_0_entry_function3,
  input  [11:0] io_decoder_0_entry_immediateOrFunction7,
  input         io_decoder_0_entry_sourceTag1_threadId,
  input  [3:0]  io_decoder_0_entry_sourceTag1_id,
  input         io_decoder_0_entry_ready1,
  input  [63:0] io_decoder_0_entry_value1,
  input         io_decoder_0_entry_sourceTag2_threadId,
  input  [3:0]  io_decoder_0_entry_sourceTag2_id,
  input         io_decoder_0_entry_ready2,
  input  [63:0] io_decoder_0_entry_value2,
  input  [3:0]  io_decoder_0_entry_destinationTag_id,
  input         io_decoder_0_entry_wasCompressed,
  input         io_decoder_0_entry_valid,
  output        io_decoder_1_ready,
  input  [6:0]  io_decoder_1_entry_opcode,
  input  [2:0]  io_decoder_1_entry_function3,
  input  [11:0] io_decoder_1_entry_immediateOrFunction7,
  input         io_decoder_1_entry_sourceTag1_threadId,
  input  [3:0]  io_decoder_1_entry_sourceTag1_id,
  input         io_decoder_1_entry_ready1,
  input  [63:0] io_decoder_1_entry_value1,
  input         io_decoder_1_entry_sourceTag2_threadId,
  input  [3:0]  io_decoder_1_entry_sourceTag2_id,
  input         io_decoder_1_entry_ready2,
  input  [63:0] io_decoder_1_entry_value2,
  input  [3:0]  io_decoder_1_entry_destinationTag_id,
  input         io_decoder_1_entry_wasCompressed,
  input         io_decoder_1_entry_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [63:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [63:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [63:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [63:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [63:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [63:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [63:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [63:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [63:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [63:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
`endif // RANDOMIZE_REG_INIT
  wire  outputArbiter_0_clock; // @[ReservationStation.scala 34:11]
  wire  outputArbiter_0_reset; // @[ReservationStation.scala 34:11]
  wire  outputArbiter_0_io_in_0_ready; // @[ReservationStation.scala 34:11]
  wire  outputArbiter_0_io_in_0_valid; // @[ReservationStation.scala 34:11]
  wire  outputArbiter_0_io_in_0_bits_destinationTag_threadId; // @[ReservationStation.scala 34:11]
  wire [3:0] outputArbiter_0_io_in_0_bits_destinationTag_id; // @[ReservationStation.scala 34:11]
  wire [63:0] outputArbiter_0_io_in_0_bits_value1; // @[ReservationStation.scala 34:11]
  wire [63:0] outputArbiter_0_io_in_0_bits_value2; // @[ReservationStation.scala 34:11]
  wire [2:0] outputArbiter_0_io_in_0_bits_function3; // @[ReservationStation.scala 34:11]
  wire [11:0] outputArbiter_0_io_in_0_bits_immediateOrFunction7; // @[ReservationStation.scala 34:11]
  wire [6:0] outputArbiter_0_io_in_0_bits_opcode; // @[ReservationStation.scala 34:11]
  wire  outputArbiter_0_io_in_0_bits_wasCompressed; // @[ReservationStation.scala 34:11]
  wire  outputArbiter_0_io_in_1_ready; // @[ReservationStation.scala 34:11]
  wire  outputArbiter_0_io_in_1_valid; // @[ReservationStation.scala 34:11]
  wire  outputArbiter_0_io_in_1_bits_destinationTag_threadId; // @[ReservationStation.scala 34:11]
  wire [3:0] outputArbiter_0_io_in_1_bits_destinationTag_id; // @[ReservationStation.scala 34:11]
  wire [63:0] outputArbiter_0_io_in_1_bits_value1; // @[ReservationStation.scala 34:11]
  wire [63:0] outputArbiter_0_io_in_1_bits_value2; // @[ReservationStation.scala 34:11]
  wire [2:0] outputArbiter_0_io_in_1_bits_function3; // @[ReservationStation.scala 34:11]
  wire [11:0] outputArbiter_0_io_in_1_bits_immediateOrFunction7; // @[ReservationStation.scala 34:11]
  wire [6:0] outputArbiter_0_io_in_1_bits_opcode; // @[ReservationStation.scala 34:11]
  wire  outputArbiter_0_io_in_1_bits_wasCompressed; // @[ReservationStation.scala 34:11]
  wire  outputArbiter_0_io_in_2_ready; // @[ReservationStation.scala 34:11]
  wire  outputArbiter_0_io_in_2_valid; // @[ReservationStation.scala 34:11]
  wire  outputArbiter_0_io_in_2_bits_destinationTag_threadId; // @[ReservationStation.scala 34:11]
  wire [3:0] outputArbiter_0_io_in_2_bits_destinationTag_id; // @[ReservationStation.scala 34:11]
  wire [63:0] outputArbiter_0_io_in_2_bits_value1; // @[ReservationStation.scala 34:11]
  wire [63:0] outputArbiter_0_io_in_2_bits_value2; // @[ReservationStation.scala 34:11]
  wire [2:0] outputArbiter_0_io_in_2_bits_function3; // @[ReservationStation.scala 34:11]
  wire [11:0] outputArbiter_0_io_in_2_bits_immediateOrFunction7; // @[ReservationStation.scala 34:11]
  wire [6:0] outputArbiter_0_io_in_2_bits_opcode; // @[ReservationStation.scala 34:11]
  wire  outputArbiter_0_io_in_2_bits_wasCompressed; // @[ReservationStation.scala 34:11]
  wire  outputArbiter_0_io_in_3_ready; // @[ReservationStation.scala 34:11]
  wire  outputArbiter_0_io_in_3_valid; // @[ReservationStation.scala 34:11]
  wire  outputArbiter_0_io_in_3_bits_destinationTag_threadId; // @[ReservationStation.scala 34:11]
  wire [3:0] outputArbiter_0_io_in_3_bits_destinationTag_id; // @[ReservationStation.scala 34:11]
  wire [63:0] outputArbiter_0_io_in_3_bits_value1; // @[ReservationStation.scala 34:11]
  wire [63:0] outputArbiter_0_io_in_3_bits_value2; // @[ReservationStation.scala 34:11]
  wire [2:0] outputArbiter_0_io_in_3_bits_function3; // @[ReservationStation.scala 34:11]
  wire [11:0] outputArbiter_0_io_in_3_bits_immediateOrFunction7; // @[ReservationStation.scala 34:11]
  wire [6:0] outputArbiter_0_io_in_3_bits_opcode; // @[ReservationStation.scala 34:11]
  wire  outputArbiter_0_io_in_3_bits_wasCompressed; // @[ReservationStation.scala 34:11]
  wire  outputArbiter_0_io_out_ready; // @[ReservationStation.scala 34:11]
  wire  outputArbiter_0_io_out_valid; // @[ReservationStation.scala 34:11]
  wire  outputArbiter_0_io_out_bits_destinationTag_threadId; // @[ReservationStation.scala 34:11]
  wire [3:0] outputArbiter_0_io_out_bits_destinationTag_id; // @[ReservationStation.scala 34:11]
  wire [63:0] outputArbiter_0_io_out_bits_value1; // @[ReservationStation.scala 34:11]
  wire [63:0] outputArbiter_0_io_out_bits_value2; // @[ReservationStation.scala 34:11]
  wire [2:0] outputArbiter_0_io_out_bits_function3; // @[ReservationStation.scala 34:11]
  wire [11:0] outputArbiter_0_io_out_bits_immediateOrFunction7; // @[ReservationStation.scala 34:11]
  wire [6:0] outputArbiter_0_io_out_bits_opcode; // @[ReservationStation.scala 34:11]
  wire  outputArbiter_0_io_out_bits_wasCompressed; // @[ReservationStation.scala 34:11]
  wire [1:0] outputArbiter_0_io_chosen; // @[ReservationStation.scala 34:11]
  wire  outputArbiter_1_clock; // @[ReservationStation.scala 34:11]
  wire  outputArbiter_1_reset; // @[ReservationStation.scala 34:11]
  wire  outputArbiter_1_io_in_0_ready; // @[ReservationStation.scala 34:11]
  wire  outputArbiter_1_io_in_0_valid; // @[ReservationStation.scala 34:11]
  wire  outputArbiter_1_io_in_0_bits_destinationTag_threadId; // @[ReservationStation.scala 34:11]
  wire [3:0] outputArbiter_1_io_in_0_bits_destinationTag_id; // @[ReservationStation.scala 34:11]
  wire [63:0] outputArbiter_1_io_in_0_bits_value1; // @[ReservationStation.scala 34:11]
  wire [63:0] outputArbiter_1_io_in_0_bits_value2; // @[ReservationStation.scala 34:11]
  wire [2:0] outputArbiter_1_io_in_0_bits_function3; // @[ReservationStation.scala 34:11]
  wire [11:0] outputArbiter_1_io_in_0_bits_immediateOrFunction7; // @[ReservationStation.scala 34:11]
  wire [6:0] outputArbiter_1_io_in_0_bits_opcode; // @[ReservationStation.scala 34:11]
  wire  outputArbiter_1_io_in_0_bits_wasCompressed; // @[ReservationStation.scala 34:11]
  wire  outputArbiter_1_io_in_1_ready; // @[ReservationStation.scala 34:11]
  wire  outputArbiter_1_io_in_1_valid; // @[ReservationStation.scala 34:11]
  wire  outputArbiter_1_io_in_1_bits_destinationTag_threadId; // @[ReservationStation.scala 34:11]
  wire [3:0] outputArbiter_1_io_in_1_bits_destinationTag_id; // @[ReservationStation.scala 34:11]
  wire [63:0] outputArbiter_1_io_in_1_bits_value1; // @[ReservationStation.scala 34:11]
  wire [63:0] outputArbiter_1_io_in_1_bits_value2; // @[ReservationStation.scala 34:11]
  wire [2:0] outputArbiter_1_io_in_1_bits_function3; // @[ReservationStation.scala 34:11]
  wire [11:0] outputArbiter_1_io_in_1_bits_immediateOrFunction7; // @[ReservationStation.scala 34:11]
  wire [6:0] outputArbiter_1_io_in_1_bits_opcode; // @[ReservationStation.scala 34:11]
  wire  outputArbiter_1_io_in_1_bits_wasCompressed; // @[ReservationStation.scala 34:11]
  wire  outputArbiter_1_io_in_2_ready; // @[ReservationStation.scala 34:11]
  wire  outputArbiter_1_io_in_2_valid; // @[ReservationStation.scala 34:11]
  wire  outputArbiter_1_io_in_2_bits_destinationTag_threadId; // @[ReservationStation.scala 34:11]
  wire [3:0] outputArbiter_1_io_in_2_bits_destinationTag_id; // @[ReservationStation.scala 34:11]
  wire [63:0] outputArbiter_1_io_in_2_bits_value1; // @[ReservationStation.scala 34:11]
  wire [63:0] outputArbiter_1_io_in_2_bits_value2; // @[ReservationStation.scala 34:11]
  wire [2:0] outputArbiter_1_io_in_2_bits_function3; // @[ReservationStation.scala 34:11]
  wire [11:0] outputArbiter_1_io_in_2_bits_immediateOrFunction7; // @[ReservationStation.scala 34:11]
  wire [6:0] outputArbiter_1_io_in_2_bits_opcode; // @[ReservationStation.scala 34:11]
  wire  outputArbiter_1_io_in_2_bits_wasCompressed; // @[ReservationStation.scala 34:11]
  wire  outputArbiter_1_io_in_3_ready; // @[ReservationStation.scala 34:11]
  wire  outputArbiter_1_io_in_3_valid; // @[ReservationStation.scala 34:11]
  wire  outputArbiter_1_io_in_3_bits_destinationTag_threadId; // @[ReservationStation.scala 34:11]
  wire [3:0] outputArbiter_1_io_in_3_bits_destinationTag_id; // @[ReservationStation.scala 34:11]
  wire [63:0] outputArbiter_1_io_in_3_bits_value1; // @[ReservationStation.scala 34:11]
  wire [63:0] outputArbiter_1_io_in_3_bits_value2; // @[ReservationStation.scala 34:11]
  wire [2:0] outputArbiter_1_io_in_3_bits_function3; // @[ReservationStation.scala 34:11]
  wire [11:0] outputArbiter_1_io_in_3_bits_immediateOrFunction7; // @[ReservationStation.scala 34:11]
  wire [6:0] outputArbiter_1_io_in_3_bits_opcode; // @[ReservationStation.scala 34:11]
  wire  outputArbiter_1_io_in_3_bits_wasCompressed; // @[ReservationStation.scala 34:11]
  wire  outputArbiter_1_io_out_ready; // @[ReservationStation.scala 34:11]
  wire  outputArbiter_1_io_out_valid; // @[ReservationStation.scala 34:11]
  wire  outputArbiter_1_io_out_bits_destinationTag_threadId; // @[ReservationStation.scala 34:11]
  wire [3:0] outputArbiter_1_io_out_bits_destinationTag_id; // @[ReservationStation.scala 34:11]
  wire [63:0] outputArbiter_1_io_out_bits_value1; // @[ReservationStation.scala 34:11]
  wire [63:0] outputArbiter_1_io_out_bits_value2; // @[ReservationStation.scala 34:11]
  wire [2:0] outputArbiter_1_io_out_bits_function3; // @[ReservationStation.scala 34:11]
  wire [11:0] outputArbiter_1_io_out_bits_immediateOrFunction7; // @[ReservationStation.scala 34:11]
  wire [6:0] outputArbiter_1_io_out_bits_opcode; // @[ReservationStation.scala 34:11]
  wire  outputArbiter_1_io_out_bits_wasCompressed; // @[ReservationStation.scala 34:11]
  wire [1:0] outputArbiter_1_io_chosen; // @[ReservationStation.scala 34:11]
  reg [6:0] reservation_0_opcode; // @[ReservationStation.scala 28:28]
  reg [2:0] reservation_0_function3; // @[ReservationStation.scala 28:28]
  reg [11:0] reservation_0_immediateOrFunction7; // @[ReservationStation.scala 28:28]
  reg  reservation_0_sourceTag1_threadId; // @[ReservationStation.scala 28:28]
  reg [3:0] reservation_0_sourceTag1_id; // @[ReservationStation.scala 28:28]
  reg  reservation_0_ready1; // @[ReservationStation.scala 28:28]
  reg [63:0] reservation_0_value1; // @[ReservationStation.scala 28:28]
  reg  reservation_0_sourceTag2_threadId; // @[ReservationStation.scala 28:28]
  reg [3:0] reservation_0_sourceTag2_id; // @[ReservationStation.scala 28:28]
  reg  reservation_0_ready2; // @[ReservationStation.scala 28:28]
  reg [63:0] reservation_0_value2; // @[ReservationStation.scala 28:28]
  reg  reservation_0_destinationTag_threadId; // @[ReservationStation.scala 28:28]
  reg [3:0] reservation_0_destinationTag_id; // @[ReservationStation.scala 28:28]
  reg  reservation_0_wasCompressed; // @[ReservationStation.scala 28:28]
  reg  reservation_0_valid; // @[ReservationStation.scala 28:28]
  reg [6:0] reservation_1_opcode; // @[ReservationStation.scala 28:28]
  reg [2:0] reservation_1_function3; // @[ReservationStation.scala 28:28]
  reg [11:0] reservation_1_immediateOrFunction7; // @[ReservationStation.scala 28:28]
  reg  reservation_1_sourceTag1_threadId; // @[ReservationStation.scala 28:28]
  reg [3:0] reservation_1_sourceTag1_id; // @[ReservationStation.scala 28:28]
  reg  reservation_1_ready1; // @[ReservationStation.scala 28:28]
  reg [63:0] reservation_1_value1; // @[ReservationStation.scala 28:28]
  reg  reservation_1_sourceTag2_threadId; // @[ReservationStation.scala 28:28]
  reg [3:0] reservation_1_sourceTag2_id; // @[ReservationStation.scala 28:28]
  reg  reservation_1_ready2; // @[ReservationStation.scala 28:28]
  reg [63:0] reservation_1_value2; // @[ReservationStation.scala 28:28]
  reg  reservation_1_destinationTag_threadId; // @[ReservationStation.scala 28:28]
  reg [3:0] reservation_1_destinationTag_id; // @[ReservationStation.scala 28:28]
  reg  reservation_1_wasCompressed; // @[ReservationStation.scala 28:28]
  reg  reservation_1_valid; // @[ReservationStation.scala 28:28]
  reg [6:0] reservation_2_opcode; // @[ReservationStation.scala 28:28]
  reg [2:0] reservation_2_function3; // @[ReservationStation.scala 28:28]
  reg [11:0] reservation_2_immediateOrFunction7; // @[ReservationStation.scala 28:28]
  reg  reservation_2_sourceTag1_threadId; // @[ReservationStation.scala 28:28]
  reg [3:0] reservation_2_sourceTag1_id; // @[ReservationStation.scala 28:28]
  reg  reservation_2_ready1; // @[ReservationStation.scala 28:28]
  reg [63:0] reservation_2_value1; // @[ReservationStation.scala 28:28]
  reg  reservation_2_sourceTag2_threadId; // @[ReservationStation.scala 28:28]
  reg [3:0] reservation_2_sourceTag2_id; // @[ReservationStation.scala 28:28]
  reg  reservation_2_ready2; // @[ReservationStation.scala 28:28]
  reg [63:0] reservation_2_value2; // @[ReservationStation.scala 28:28]
  reg  reservation_2_destinationTag_threadId; // @[ReservationStation.scala 28:28]
  reg [3:0] reservation_2_destinationTag_id; // @[ReservationStation.scala 28:28]
  reg  reservation_2_wasCompressed; // @[ReservationStation.scala 28:28]
  reg  reservation_2_valid; // @[ReservationStation.scala 28:28]
  reg [6:0] reservation_3_opcode; // @[ReservationStation.scala 28:28]
  reg [2:0] reservation_3_function3; // @[ReservationStation.scala 28:28]
  reg [11:0] reservation_3_immediateOrFunction7; // @[ReservationStation.scala 28:28]
  reg  reservation_3_sourceTag1_threadId; // @[ReservationStation.scala 28:28]
  reg [3:0] reservation_3_sourceTag1_id; // @[ReservationStation.scala 28:28]
  reg  reservation_3_ready1; // @[ReservationStation.scala 28:28]
  reg [63:0] reservation_3_value1; // @[ReservationStation.scala 28:28]
  reg  reservation_3_sourceTag2_threadId; // @[ReservationStation.scala 28:28]
  reg [3:0] reservation_3_sourceTag2_id; // @[ReservationStation.scala 28:28]
  reg  reservation_3_ready2; // @[ReservationStation.scala 28:28]
  reg [63:0] reservation_3_value2; // @[ReservationStation.scala 28:28]
  reg  reservation_3_destinationTag_threadId; // @[ReservationStation.scala 28:28]
  reg [3:0] reservation_3_destinationTag_id; // @[ReservationStation.scala 28:28]
  reg  reservation_3_wasCompressed; // @[ReservationStation.scala 28:28]
  reg  reservation_3_valid; // @[ReservationStation.scala 28:28]
  reg [6:0] reservation_4_opcode; // @[ReservationStation.scala 28:28]
  reg [2:0] reservation_4_function3; // @[ReservationStation.scala 28:28]
  reg [11:0] reservation_4_immediateOrFunction7; // @[ReservationStation.scala 28:28]
  reg  reservation_4_sourceTag1_threadId; // @[ReservationStation.scala 28:28]
  reg [3:0] reservation_4_sourceTag1_id; // @[ReservationStation.scala 28:28]
  reg  reservation_4_ready1; // @[ReservationStation.scala 28:28]
  reg [63:0] reservation_4_value1; // @[ReservationStation.scala 28:28]
  reg  reservation_4_sourceTag2_threadId; // @[ReservationStation.scala 28:28]
  reg [3:0] reservation_4_sourceTag2_id; // @[ReservationStation.scala 28:28]
  reg  reservation_4_ready2; // @[ReservationStation.scala 28:28]
  reg [63:0] reservation_4_value2; // @[ReservationStation.scala 28:28]
  reg  reservation_4_destinationTag_threadId; // @[ReservationStation.scala 28:28]
  reg [3:0] reservation_4_destinationTag_id; // @[ReservationStation.scala 28:28]
  reg  reservation_4_wasCompressed; // @[ReservationStation.scala 28:28]
  reg  reservation_4_valid; // @[ReservationStation.scala 28:28]
  reg [6:0] reservation_5_opcode; // @[ReservationStation.scala 28:28]
  reg [2:0] reservation_5_function3; // @[ReservationStation.scala 28:28]
  reg [11:0] reservation_5_immediateOrFunction7; // @[ReservationStation.scala 28:28]
  reg  reservation_5_sourceTag1_threadId; // @[ReservationStation.scala 28:28]
  reg [3:0] reservation_5_sourceTag1_id; // @[ReservationStation.scala 28:28]
  reg  reservation_5_ready1; // @[ReservationStation.scala 28:28]
  reg [63:0] reservation_5_value1; // @[ReservationStation.scala 28:28]
  reg  reservation_5_sourceTag2_threadId; // @[ReservationStation.scala 28:28]
  reg [3:0] reservation_5_sourceTag2_id; // @[ReservationStation.scala 28:28]
  reg  reservation_5_ready2; // @[ReservationStation.scala 28:28]
  reg [63:0] reservation_5_value2; // @[ReservationStation.scala 28:28]
  reg  reservation_5_destinationTag_threadId; // @[ReservationStation.scala 28:28]
  reg [3:0] reservation_5_destinationTag_id; // @[ReservationStation.scala 28:28]
  reg  reservation_5_wasCompressed; // @[ReservationStation.scala 28:28]
  reg  reservation_5_valid; // @[ReservationStation.scala 28:28]
  reg [6:0] reservation_6_opcode; // @[ReservationStation.scala 28:28]
  reg [2:0] reservation_6_function3; // @[ReservationStation.scala 28:28]
  reg [11:0] reservation_6_immediateOrFunction7; // @[ReservationStation.scala 28:28]
  reg  reservation_6_sourceTag1_threadId; // @[ReservationStation.scala 28:28]
  reg [3:0] reservation_6_sourceTag1_id; // @[ReservationStation.scala 28:28]
  reg  reservation_6_ready1; // @[ReservationStation.scala 28:28]
  reg [63:0] reservation_6_value1; // @[ReservationStation.scala 28:28]
  reg  reservation_6_sourceTag2_threadId; // @[ReservationStation.scala 28:28]
  reg [3:0] reservation_6_sourceTag2_id; // @[ReservationStation.scala 28:28]
  reg  reservation_6_ready2; // @[ReservationStation.scala 28:28]
  reg [63:0] reservation_6_value2; // @[ReservationStation.scala 28:28]
  reg  reservation_6_destinationTag_threadId; // @[ReservationStation.scala 28:28]
  reg [3:0] reservation_6_destinationTag_id; // @[ReservationStation.scala 28:28]
  reg  reservation_6_wasCompressed; // @[ReservationStation.scala 28:28]
  reg  reservation_6_valid; // @[ReservationStation.scala 28:28]
  reg [6:0] reservation_7_opcode; // @[ReservationStation.scala 28:28]
  reg [2:0] reservation_7_function3; // @[ReservationStation.scala 28:28]
  reg [11:0] reservation_7_immediateOrFunction7; // @[ReservationStation.scala 28:28]
  reg  reservation_7_sourceTag1_threadId; // @[ReservationStation.scala 28:28]
  reg [3:0] reservation_7_sourceTag1_id; // @[ReservationStation.scala 28:28]
  reg  reservation_7_ready1; // @[ReservationStation.scala 28:28]
  reg [63:0] reservation_7_value1; // @[ReservationStation.scala 28:28]
  reg  reservation_7_sourceTag2_threadId; // @[ReservationStation.scala 28:28]
  reg [3:0] reservation_7_sourceTag2_id; // @[ReservationStation.scala 28:28]
  reg  reservation_7_ready2; // @[ReservationStation.scala 28:28]
  reg [63:0] reservation_7_value2; // @[ReservationStation.scala 28:28]
  reg  reservation_7_destinationTag_threadId; // @[ReservationStation.scala 28:28]
  reg [3:0] reservation_7_destinationTag_id; // @[ReservationStation.scala 28:28]
  reg  reservation_7_wasCompressed; // @[ReservationStation.scala 28:28]
  reg  reservation_7_valid; // @[ReservationStation.scala 28:28]
  wire  _GEN_0 = outputArbiter_0_io_in_0_valid & outputArbiter_0_io_in_0_ready ? 1'h0 : reservation_0_valid; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire  _GEN_1 = outputArbiter_0_io_in_0_valid & outputArbiter_0_io_in_0_ready ? 1'h0 : reservation_0_wasCompressed; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire [3:0] _GEN_2 = outputArbiter_0_io_in_0_valid & outputArbiter_0_io_in_0_ready ? 4'h0 :
    reservation_0_destinationTag_id; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire  _GEN_3 = outputArbiter_0_io_in_0_valid & outputArbiter_0_io_in_0_ready ? 1'h0 :
    reservation_0_destinationTag_threadId; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire [63:0] _GEN_4 = outputArbiter_0_io_in_0_valid & outputArbiter_0_io_in_0_ready ? 64'h0 : reservation_0_value2; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire  _GEN_5 = outputArbiter_0_io_in_0_valid & outputArbiter_0_io_in_0_ready ? 1'h0 : reservation_0_ready2; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire [3:0] _GEN_6 = outputArbiter_0_io_in_0_valid & outputArbiter_0_io_in_0_ready ? 4'h0 : reservation_0_sourceTag2_id
    ; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire  _GEN_7 = outputArbiter_0_io_in_0_valid & outputArbiter_0_io_in_0_ready ? 1'h0 :
    reservation_0_sourceTag2_threadId; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire [63:0] _GEN_8 = outputArbiter_0_io_in_0_valid & outputArbiter_0_io_in_0_ready ? 64'h0 : reservation_0_value1; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire  _GEN_9 = outputArbiter_0_io_in_0_valid & outputArbiter_0_io_in_0_ready ? 1'h0 : reservation_0_ready1; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire [3:0] _GEN_10 = outputArbiter_0_io_in_0_valid & outputArbiter_0_io_in_0_ready ? 4'h0 :
    reservation_0_sourceTag1_id; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire  _GEN_11 = outputArbiter_0_io_in_0_valid & outputArbiter_0_io_in_0_ready ? 1'h0 :
    reservation_0_sourceTag1_threadId; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire [11:0] _GEN_12 = outputArbiter_0_io_in_0_valid & outputArbiter_0_io_in_0_ready ? 12'h0 :
    reservation_0_immediateOrFunction7; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire [2:0] _GEN_13 = outputArbiter_0_io_in_0_valid & outputArbiter_0_io_in_0_ready ? 3'h0 : reservation_0_function3; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire [6:0] _GEN_14 = outputArbiter_0_io_in_0_valid & outputArbiter_0_io_in_0_ready ? 7'h0 : reservation_0_opcode; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire  _GEN_15 = outputArbiter_0_io_in_1_valid & outputArbiter_0_io_in_1_ready ? 1'h0 : reservation_2_valid; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire  _GEN_16 = outputArbiter_0_io_in_1_valid & outputArbiter_0_io_in_1_ready ? 1'h0 : reservation_2_wasCompressed; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire [3:0] _GEN_17 = outputArbiter_0_io_in_1_valid & outputArbiter_0_io_in_1_ready ? 4'h0 :
    reservation_2_destinationTag_id; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire  _GEN_18 = outputArbiter_0_io_in_1_valid & outputArbiter_0_io_in_1_ready ? 1'h0 :
    reservation_2_destinationTag_threadId; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire [63:0] _GEN_19 = outputArbiter_0_io_in_1_valid & outputArbiter_0_io_in_1_ready ? 64'h0 : reservation_2_value2; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire  _GEN_20 = outputArbiter_0_io_in_1_valid & outputArbiter_0_io_in_1_ready ? 1'h0 : reservation_2_ready2; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire [3:0] _GEN_21 = outputArbiter_0_io_in_1_valid & outputArbiter_0_io_in_1_ready ? 4'h0 :
    reservation_2_sourceTag2_id; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire  _GEN_22 = outputArbiter_0_io_in_1_valid & outputArbiter_0_io_in_1_ready ? 1'h0 :
    reservation_2_sourceTag2_threadId; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire [63:0] _GEN_23 = outputArbiter_0_io_in_1_valid & outputArbiter_0_io_in_1_ready ? 64'h0 : reservation_2_value1; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire  _GEN_24 = outputArbiter_0_io_in_1_valid & outputArbiter_0_io_in_1_ready ? 1'h0 : reservation_2_ready1; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire [3:0] _GEN_25 = outputArbiter_0_io_in_1_valid & outputArbiter_0_io_in_1_ready ? 4'h0 :
    reservation_2_sourceTag1_id; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire  _GEN_26 = outputArbiter_0_io_in_1_valid & outputArbiter_0_io_in_1_ready ? 1'h0 :
    reservation_2_sourceTag1_threadId; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire [11:0] _GEN_27 = outputArbiter_0_io_in_1_valid & outputArbiter_0_io_in_1_ready ? 12'h0 :
    reservation_2_immediateOrFunction7; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire [2:0] _GEN_28 = outputArbiter_0_io_in_1_valid & outputArbiter_0_io_in_1_ready ? 3'h0 : reservation_2_function3; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire [6:0] _GEN_29 = outputArbiter_0_io_in_1_valid & outputArbiter_0_io_in_1_ready ? 7'h0 : reservation_2_opcode; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire  _GEN_30 = outputArbiter_0_io_in_2_valid & outputArbiter_0_io_in_2_ready ? 1'h0 : reservation_4_valid; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire  _GEN_31 = outputArbiter_0_io_in_2_valid & outputArbiter_0_io_in_2_ready ? 1'h0 : reservation_4_wasCompressed; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire [3:0] _GEN_32 = outputArbiter_0_io_in_2_valid & outputArbiter_0_io_in_2_ready ? 4'h0 :
    reservation_4_destinationTag_id; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire  _GEN_33 = outputArbiter_0_io_in_2_valid & outputArbiter_0_io_in_2_ready ? 1'h0 :
    reservation_4_destinationTag_threadId; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire [63:0] _GEN_34 = outputArbiter_0_io_in_2_valid & outputArbiter_0_io_in_2_ready ? 64'h0 : reservation_4_value2; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire  _GEN_35 = outputArbiter_0_io_in_2_valid & outputArbiter_0_io_in_2_ready ? 1'h0 : reservation_4_ready2; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire [3:0] _GEN_36 = outputArbiter_0_io_in_2_valid & outputArbiter_0_io_in_2_ready ? 4'h0 :
    reservation_4_sourceTag2_id; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire  _GEN_37 = outputArbiter_0_io_in_2_valid & outputArbiter_0_io_in_2_ready ? 1'h0 :
    reservation_4_sourceTag2_threadId; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire [63:0] _GEN_38 = outputArbiter_0_io_in_2_valid & outputArbiter_0_io_in_2_ready ? 64'h0 : reservation_4_value1; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire  _GEN_39 = outputArbiter_0_io_in_2_valid & outputArbiter_0_io_in_2_ready ? 1'h0 : reservation_4_ready1; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire [3:0] _GEN_40 = outputArbiter_0_io_in_2_valid & outputArbiter_0_io_in_2_ready ? 4'h0 :
    reservation_4_sourceTag1_id; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire  _GEN_41 = outputArbiter_0_io_in_2_valid & outputArbiter_0_io_in_2_ready ? 1'h0 :
    reservation_4_sourceTag1_threadId; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire [11:0] _GEN_42 = outputArbiter_0_io_in_2_valid & outputArbiter_0_io_in_2_ready ? 12'h0 :
    reservation_4_immediateOrFunction7; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire [2:0] _GEN_43 = outputArbiter_0_io_in_2_valid & outputArbiter_0_io_in_2_ready ? 3'h0 : reservation_4_function3; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire [6:0] _GEN_44 = outputArbiter_0_io_in_2_valid & outputArbiter_0_io_in_2_ready ? 7'h0 : reservation_4_opcode; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire  _GEN_45 = outputArbiter_0_io_in_3_valid & outputArbiter_0_io_in_3_ready ? 1'h0 : reservation_6_valid; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire  _GEN_46 = outputArbiter_0_io_in_3_valid & outputArbiter_0_io_in_3_ready ? 1'h0 : reservation_6_wasCompressed; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire [3:0] _GEN_47 = outputArbiter_0_io_in_3_valid & outputArbiter_0_io_in_3_ready ? 4'h0 :
    reservation_6_destinationTag_id; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire  _GEN_48 = outputArbiter_0_io_in_3_valid & outputArbiter_0_io_in_3_ready ? 1'h0 :
    reservation_6_destinationTag_threadId; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire [63:0] _GEN_49 = outputArbiter_0_io_in_3_valid & outputArbiter_0_io_in_3_ready ? 64'h0 : reservation_6_value2; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire  _GEN_50 = outputArbiter_0_io_in_3_valid & outputArbiter_0_io_in_3_ready ? 1'h0 : reservation_6_ready2; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire [3:0] _GEN_51 = outputArbiter_0_io_in_3_valid & outputArbiter_0_io_in_3_ready ? 4'h0 :
    reservation_6_sourceTag2_id; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire  _GEN_52 = outputArbiter_0_io_in_3_valid & outputArbiter_0_io_in_3_ready ? 1'h0 :
    reservation_6_sourceTag2_threadId; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire [63:0] _GEN_53 = outputArbiter_0_io_in_3_valid & outputArbiter_0_io_in_3_ready ? 64'h0 : reservation_6_value1; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire  _GEN_54 = outputArbiter_0_io_in_3_valid & outputArbiter_0_io_in_3_ready ? 1'h0 : reservation_6_ready1; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire [3:0] _GEN_55 = outputArbiter_0_io_in_3_valid & outputArbiter_0_io_in_3_ready ? 4'h0 :
    reservation_6_sourceTag1_id; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire  _GEN_56 = outputArbiter_0_io_in_3_valid & outputArbiter_0_io_in_3_ready ? 1'h0 :
    reservation_6_sourceTag1_threadId; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire [11:0] _GEN_57 = outputArbiter_0_io_in_3_valid & outputArbiter_0_io_in_3_ready ? 12'h0 :
    reservation_6_immediateOrFunction7; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire [2:0] _GEN_58 = outputArbiter_0_io_in_3_valid & outputArbiter_0_io_in_3_ready ? 3'h0 : reservation_6_function3; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire [6:0] _GEN_59 = outputArbiter_0_io_in_3_valid & outputArbiter_0_io_in_3_ready ? 7'h0 : reservation_6_opcode; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire  _GEN_60 = outputArbiter_1_io_in_0_valid & outputArbiter_1_io_in_0_ready ? 1'h0 : reservation_1_valid; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire  _GEN_61 = outputArbiter_1_io_in_0_valid & outputArbiter_1_io_in_0_ready ? 1'h0 : reservation_1_wasCompressed; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire [3:0] _GEN_62 = outputArbiter_1_io_in_0_valid & outputArbiter_1_io_in_0_ready ? 4'h0 :
    reservation_1_destinationTag_id; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire  _GEN_63 = outputArbiter_1_io_in_0_valid & outputArbiter_1_io_in_0_ready ? 1'h0 :
    reservation_1_destinationTag_threadId; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire [63:0] _GEN_64 = outputArbiter_1_io_in_0_valid & outputArbiter_1_io_in_0_ready ? 64'h0 : reservation_1_value2; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire  _GEN_65 = outputArbiter_1_io_in_0_valid & outputArbiter_1_io_in_0_ready ? 1'h0 : reservation_1_ready2; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire [3:0] _GEN_66 = outputArbiter_1_io_in_0_valid & outputArbiter_1_io_in_0_ready ? 4'h0 :
    reservation_1_sourceTag2_id; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire  _GEN_67 = outputArbiter_1_io_in_0_valid & outputArbiter_1_io_in_0_ready ? 1'h0 :
    reservation_1_sourceTag2_threadId; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire [63:0] _GEN_68 = outputArbiter_1_io_in_0_valid & outputArbiter_1_io_in_0_ready ? 64'h0 : reservation_1_value1; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire  _GEN_69 = outputArbiter_1_io_in_0_valid & outputArbiter_1_io_in_0_ready ? 1'h0 : reservation_1_ready1; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire [3:0] _GEN_70 = outputArbiter_1_io_in_0_valid & outputArbiter_1_io_in_0_ready ? 4'h0 :
    reservation_1_sourceTag1_id; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire  _GEN_71 = outputArbiter_1_io_in_0_valid & outputArbiter_1_io_in_0_ready ? 1'h0 :
    reservation_1_sourceTag1_threadId; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire [11:0] _GEN_72 = outputArbiter_1_io_in_0_valid & outputArbiter_1_io_in_0_ready ? 12'h0 :
    reservation_1_immediateOrFunction7; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire [2:0] _GEN_73 = outputArbiter_1_io_in_0_valid & outputArbiter_1_io_in_0_ready ? 3'h0 : reservation_1_function3; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire [6:0] _GEN_74 = outputArbiter_1_io_in_0_valid & outputArbiter_1_io_in_0_ready ? 7'h0 : reservation_1_opcode; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire  _GEN_75 = outputArbiter_1_io_in_1_valid & outputArbiter_1_io_in_1_ready ? 1'h0 : reservation_3_valid; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire  _GEN_76 = outputArbiter_1_io_in_1_valid & outputArbiter_1_io_in_1_ready ? 1'h0 : reservation_3_wasCompressed; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire [3:0] _GEN_77 = outputArbiter_1_io_in_1_valid & outputArbiter_1_io_in_1_ready ? 4'h0 :
    reservation_3_destinationTag_id; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire  _GEN_78 = outputArbiter_1_io_in_1_valid & outputArbiter_1_io_in_1_ready ? 1'h0 :
    reservation_3_destinationTag_threadId; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire [63:0] _GEN_79 = outputArbiter_1_io_in_1_valid & outputArbiter_1_io_in_1_ready ? 64'h0 : reservation_3_value2; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire  _GEN_80 = outputArbiter_1_io_in_1_valid & outputArbiter_1_io_in_1_ready ? 1'h0 : reservation_3_ready2; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire [3:0] _GEN_81 = outputArbiter_1_io_in_1_valid & outputArbiter_1_io_in_1_ready ? 4'h0 :
    reservation_3_sourceTag2_id; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire  _GEN_82 = outputArbiter_1_io_in_1_valid & outputArbiter_1_io_in_1_ready ? 1'h0 :
    reservation_3_sourceTag2_threadId; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire [63:0] _GEN_83 = outputArbiter_1_io_in_1_valid & outputArbiter_1_io_in_1_ready ? 64'h0 : reservation_3_value1; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire  _GEN_84 = outputArbiter_1_io_in_1_valid & outputArbiter_1_io_in_1_ready ? 1'h0 : reservation_3_ready1; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire [3:0] _GEN_85 = outputArbiter_1_io_in_1_valid & outputArbiter_1_io_in_1_ready ? 4'h0 :
    reservation_3_sourceTag1_id; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire  _GEN_86 = outputArbiter_1_io_in_1_valid & outputArbiter_1_io_in_1_ready ? 1'h0 :
    reservation_3_sourceTag1_threadId; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire [11:0] _GEN_87 = outputArbiter_1_io_in_1_valid & outputArbiter_1_io_in_1_ready ? 12'h0 :
    reservation_3_immediateOrFunction7; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire [2:0] _GEN_88 = outputArbiter_1_io_in_1_valid & outputArbiter_1_io_in_1_ready ? 3'h0 : reservation_3_function3; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire [6:0] _GEN_89 = outputArbiter_1_io_in_1_valid & outputArbiter_1_io_in_1_ready ? 7'h0 : reservation_3_opcode; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire  _GEN_90 = outputArbiter_1_io_in_2_valid & outputArbiter_1_io_in_2_ready ? 1'h0 : reservation_5_valid; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire  _GEN_91 = outputArbiter_1_io_in_2_valid & outputArbiter_1_io_in_2_ready ? 1'h0 : reservation_5_wasCompressed; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire [3:0] _GEN_92 = outputArbiter_1_io_in_2_valid & outputArbiter_1_io_in_2_ready ? 4'h0 :
    reservation_5_destinationTag_id; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire  _GEN_93 = outputArbiter_1_io_in_2_valid & outputArbiter_1_io_in_2_ready ? 1'h0 :
    reservation_5_destinationTag_threadId; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire [63:0] _GEN_94 = outputArbiter_1_io_in_2_valid & outputArbiter_1_io_in_2_ready ? 64'h0 : reservation_5_value2; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire  _GEN_95 = outputArbiter_1_io_in_2_valid & outputArbiter_1_io_in_2_ready ? 1'h0 : reservation_5_ready2; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire [3:0] _GEN_96 = outputArbiter_1_io_in_2_valid & outputArbiter_1_io_in_2_ready ? 4'h0 :
    reservation_5_sourceTag2_id; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire  _GEN_97 = outputArbiter_1_io_in_2_valid & outputArbiter_1_io_in_2_ready ? 1'h0 :
    reservation_5_sourceTag2_threadId; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire [63:0] _GEN_98 = outputArbiter_1_io_in_2_valid & outputArbiter_1_io_in_2_ready ? 64'h0 : reservation_5_value1; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire  _GEN_99 = outputArbiter_1_io_in_2_valid & outputArbiter_1_io_in_2_ready ? 1'h0 : reservation_5_ready1; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire [3:0] _GEN_100 = outputArbiter_1_io_in_2_valid & outputArbiter_1_io_in_2_ready ? 4'h0 :
    reservation_5_sourceTag1_id; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire  _GEN_101 = outputArbiter_1_io_in_2_valid & outputArbiter_1_io_in_2_ready ? 1'h0 :
    reservation_5_sourceTag1_threadId; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire [11:0] _GEN_102 = outputArbiter_1_io_in_2_valid & outputArbiter_1_io_in_2_ready ? 12'h0 :
    reservation_5_immediateOrFunction7; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire [2:0] _GEN_103 = outputArbiter_1_io_in_2_valid & outputArbiter_1_io_in_2_ready ? 3'h0 : reservation_5_function3; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire [6:0] _GEN_104 = outputArbiter_1_io_in_2_valid & outputArbiter_1_io_in_2_ready ? 7'h0 : reservation_5_opcode; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire  _GEN_105 = outputArbiter_1_io_in_3_valid & outputArbiter_1_io_in_3_ready ? 1'h0 : reservation_7_valid; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire  _GEN_106 = outputArbiter_1_io_in_3_valid & outputArbiter_1_io_in_3_ready ? 1'h0 : reservation_7_wasCompressed; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire [3:0] _GEN_107 = outputArbiter_1_io_in_3_valid & outputArbiter_1_io_in_3_ready ? 4'h0 :
    reservation_7_destinationTag_id; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire  _GEN_108 = outputArbiter_1_io_in_3_valid & outputArbiter_1_io_in_3_ready ? 1'h0 :
    reservation_7_destinationTag_threadId; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire [63:0] _GEN_109 = outputArbiter_1_io_in_3_valid & outputArbiter_1_io_in_3_ready ? 64'h0 : reservation_7_value2; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire  _GEN_110 = outputArbiter_1_io_in_3_valid & outputArbiter_1_io_in_3_ready ? 1'h0 : reservation_7_ready2; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire [3:0] _GEN_111 = outputArbiter_1_io_in_3_valid & outputArbiter_1_io_in_3_ready ? 4'h0 :
    reservation_7_sourceTag2_id; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire  _GEN_112 = outputArbiter_1_io_in_3_valid & outputArbiter_1_io_in_3_ready ? 1'h0 :
    reservation_7_sourceTag2_threadId; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire [63:0] _GEN_113 = outputArbiter_1_io_in_3_valid & outputArbiter_1_io_in_3_ready ? 64'h0 : reservation_7_value1; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire  _GEN_114 = outputArbiter_1_io_in_3_valid & outputArbiter_1_io_in_3_ready ? 1'h0 : reservation_7_ready1; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire [3:0] _GEN_115 = outputArbiter_1_io_in_3_valid & outputArbiter_1_io_in_3_ready ? 4'h0 :
    reservation_7_sourceTag1_id; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire  _GEN_116 = outputArbiter_1_io_in_3_valid & outputArbiter_1_io_in_3_ready ? 1'h0 :
    reservation_7_sourceTag1_threadId; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire [11:0] _GEN_117 = outputArbiter_1_io_in_3_valid & outputArbiter_1_io_in_3_ready ? 12'h0 :
    reservation_7_immediateOrFunction7; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire [2:0] _GEN_118 = outputArbiter_1_io_in_3_valid & outputArbiter_1_io_in_3_ready ? 3'h0 : reservation_7_function3; // @[ReservationStation.scala 54:32 55:11 28:28]
  wire [6:0] _GEN_119 = outputArbiter_1_io_in_3_valid & outputArbiter_1_io_in_3_ready ? 7'h0 : reservation_7_opcode; // @[ReservationStation.scala 54:32 55:11 28:28]
  reg [2:0] head; // @[ReservationStation.scala 62:29]
  wire  _GEN_121 = 3'h1 == head ? reservation_1_valid : reservation_0_valid; // @[ReservationStation.scala 66:{10,10}]
  wire  _GEN_122 = 3'h2 == head ? reservation_2_valid : _GEN_121; // @[ReservationStation.scala 66:{10,10}]
  wire  _GEN_123 = 3'h3 == head ? reservation_3_valid : _GEN_122; // @[ReservationStation.scala 66:{10,10}]
  wire  _GEN_124 = 3'h4 == head ? reservation_4_valid : _GEN_123; // @[ReservationStation.scala 66:{10,10}]
  wire  _GEN_125 = 3'h5 == head ? reservation_5_valid : _GEN_124; // @[ReservationStation.scala 66:{10,10}]
  wire  _GEN_126 = 3'h6 == head ? reservation_6_valid : _GEN_125; // @[ReservationStation.scala 66:{10,10}]
  wire  _GEN_127 = 3'h7 == head ? reservation_7_valid : _GEN_126; // @[ReservationStation.scala 66:{10,10}]
  wire  _T_8 = ~_GEN_127; // @[ReservationStation.scala 66:10]
  wire [6:0] _GEN_128 = 3'h0 == head ? io_decoder_0_entry_opcode : _GEN_14; // @[ReservationStation.scala 69:{31,31}]
  wire [6:0] _GEN_129 = 3'h1 == head ? io_decoder_0_entry_opcode : _GEN_74; // @[ReservationStation.scala 69:{31,31}]
  wire [6:0] _GEN_130 = 3'h2 == head ? io_decoder_0_entry_opcode : _GEN_29; // @[ReservationStation.scala 69:{31,31}]
  wire [6:0] _GEN_131 = 3'h3 == head ? io_decoder_0_entry_opcode : _GEN_89; // @[ReservationStation.scala 69:{31,31}]
  wire [6:0] _GEN_132 = 3'h4 == head ? io_decoder_0_entry_opcode : _GEN_44; // @[ReservationStation.scala 69:{31,31}]
  wire [6:0] _GEN_133 = 3'h5 == head ? io_decoder_0_entry_opcode : _GEN_104; // @[ReservationStation.scala 69:{31,31}]
  wire [6:0] _GEN_134 = 3'h6 == head ? io_decoder_0_entry_opcode : _GEN_59; // @[ReservationStation.scala 69:{31,31}]
  wire [6:0] _GEN_135 = 3'h7 == head ? io_decoder_0_entry_opcode : _GEN_119; // @[ReservationStation.scala 69:{31,31}]
  wire [2:0] _GEN_136 = 3'h0 == head ? io_decoder_0_entry_function3 : _GEN_13; // @[ReservationStation.scala 69:{31,31}]
  wire [2:0] _GEN_137 = 3'h1 == head ? io_decoder_0_entry_function3 : _GEN_73; // @[ReservationStation.scala 69:{31,31}]
  wire [2:0] _GEN_138 = 3'h2 == head ? io_decoder_0_entry_function3 : _GEN_28; // @[ReservationStation.scala 69:{31,31}]
  wire [2:0] _GEN_139 = 3'h3 == head ? io_decoder_0_entry_function3 : _GEN_88; // @[ReservationStation.scala 69:{31,31}]
  wire [2:0] _GEN_140 = 3'h4 == head ? io_decoder_0_entry_function3 : _GEN_43; // @[ReservationStation.scala 69:{31,31}]
  wire [2:0] _GEN_141 = 3'h5 == head ? io_decoder_0_entry_function3 : _GEN_103; // @[ReservationStation.scala 69:{31,31}]
  wire [2:0] _GEN_142 = 3'h6 == head ? io_decoder_0_entry_function3 : _GEN_58; // @[ReservationStation.scala 69:{31,31}]
  wire [2:0] _GEN_143 = 3'h7 == head ? io_decoder_0_entry_function3 : _GEN_118; // @[ReservationStation.scala 69:{31,31}]
  wire [11:0] _GEN_144 = 3'h0 == head ? io_decoder_0_entry_immediateOrFunction7 : _GEN_12; // @[ReservationStation.scala 69:{31,31}]
  wire [11:0] _GEN_145 = 3'h1 == head ? io_decoder_0_entry_immediateOrFunction7 : _GEN_72; // @[ReservationStation.scala 69:{31,31}]
  wire [11:0] _GEN_146 = 3'h2 == head ? io_decoder_0_entry_immediateOrFunction7 : _GEN_27; // @[ReservationStation.scala 69:{31,31}]
  wire [11:0] _GEN_147 = 3'h3 == head ? io_decoder_0_entry_immediateOrFunction7 : _GEN_87; // @[ReservationStation.scala 69:{31,31}]
  wire [11:0] _GEN_148 = 3'h4 == head ? io_decoder_0_entry_immediateOrFunction7 : _GEN_42; // @[ReservationStation.scala 69:{31,31}]
  wire [11:0] _GEN_149 = 3'h5 == head ? io_decoder_0_entry_immediateOrFunction7 : _GEN_102; // @[ReservationStation.scala 69:{31,31}]
  wire [11:0] _GEN_150 = 3'h6 == head ? io_decoder_0_entry_immediateOrFunction7 : _GEN_57; // @[ReservationStation.scala 69:{31,31}]
  wire [11:0] _GEN_151 = 3'h7 == head ? io_decoder_0_entry_immediateOrFunction7 : _GEN_117; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_152 = 3'h0 == head ? io_decoder_0_entry_sourceTag1_threadId : _GEN_11; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_153 = 3'h1 == head ? io_decoder_0_entry_sourceTag1_threadId : _GEN_71; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_154 = 3'h2 == head ? io_decoder_0_entry_sourceTag1_threadId : _GEN_26; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_155 = 3'h3 == head ? io_decoder_0_entry_sourceTag1_threadId : _GEN_86; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_156 = 3'h4 == head ? io_decoder_0_entry_sourceTag1_threadId : _GEN_41; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_157 = 3'h5 == head ? io_decoder_0_entry_sourceTag1_threadId : _GEN_101; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_158 = 3'h6 == head ? io_decoder_0_entry_sourceTag1_threadId : _GEN_56; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_159 = 3'h7 == head ? io_decoder_0_entry_sourceTag1_threadId : _GEN_116; // @[ReservationStation.scala 69:{31,31}]
  wire [3:0] _GEN_160 = 3'h0 == head ? io_decoder_0_entry_sourceTag1_id : _GEN_10; // @[ReservationStation.scala 69:{31,31}]
  wire [3:0] _GEN_161 = 3'h1 == head ? io_decoder_0_entry_sourceTag1_id : _GEN_70; // @[ReservationStation.scala 69:{31,31}]
  wire [3:0] _GEN_162 = 3'h2 == head ? io_decoder_0_entry_sourceTag1_id : _GEN_25; // @[ReservationStation.scala 69:{31,31}]
  wire [3:0] _GEN_163 = 3'h3 == head ? io_decoder_0_entry_sourceTag1_id : _GEN_85; // @[ReservationStation.scala 69:{31,31}]
  wire [3:0] _GEN_164 = 3'h4 == head ? io_decoder_0_entry_sourceTag1_id : _GEN_40; // @[ReservationStation.scala 69:{31,31}]
  wire [3:0] _GEN_165 = 3'h5 == head ? io_decoder_0_entry_sourceTag1_id : _GEN_100; // @[ReservationStation.scala 69:{31,31}]
  wire [3:0] _GEN_166 = 3'h6 == head ? io_decoder_0_entry_sourceTag1_id : _GEN_55; // @[ReservationStation.scala 69:{31,31}]
  wire [3:0] _GEN_167 = 3'h7 == head ? io_decoder_0_entry_sourceTag1_id : _GEN_115; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_168 = 3'h0 == head ? io_decoder_0_entry_ready1 : _GEN_9; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_169 = 3'h1 == head ? io_decoder_0_entry_ready1 : _GEN_69; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_170 = 3'h2 == head ? io_decoder_0_entry_ready1 : _GEN_24; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_171 = 3'h3 == head ? io_decoder_0_entry_ready1 : _GEN_84; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_172 = 3'h4 == head ? io_decoder_0_entry_ready1 : _GEN_39; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_173 = 3'h5 == head ? io_decoder_0_entry_ready1 : _GEN_99; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_174 = 3'h6 == head ? io_decoder_0_entry_ready1 : _GEN_54; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_175 = 3'h7 == head ? io_decoder_0_entry_ready1 : _GEN_114; // @[ReservationStation.scala 69:{31,31}]
  wire [63:0] _GEN_176 = 3'h0 == head ? io_decoder_0_entry_value1 : _GEN_8; // @[ReservationStation.scala 69:{31,31}]
  wire [63:0] _GEN_177 = 3'h1 == head ? io_decoder_0_entry_value1 : _GEN_68; // @[ReservationStation.scala 69:{31,31}]
  wire [63:0] _GEN_178 = 3'h2 == head ? io_decoder_0_entry_value1 : _GEN_23; // @[ReservationStation.scala 69:{31,31}]
  wire [63:0] _GEN_179 = 3'h3 == head ? io_decoder_0_entry_value1 : _GEN_83; // @[ReservationStation.scala 69:{31,31}]
  wire [63:0] _GEN_180 = 3'h4 == head ? io_decoder_0_entry_value1 : _GEN_38; // @[ReservationStation.scala 69:{31,31}]
  wire [63:0] _GEN_181 = 3'h5 == head ? io_decoder_0_entry_value1 : _GEN_98; // @[ReservationStation.scala 69:{31,31}]
  wire [63:0] _GEN_182 = 3'h6 == head ? io_decoder_0_entry_value1 : _GEN_53; // @[ReservationStation.scala 69:{31,31}]
  wire [63:0] _GEN_183 = 3'h7 == head ? io_decoder_0_entry_value1 : _GEN_113; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_184 = 3'h0 == head ? io_decoder_0_entry_sourceTag2_threadId : _GEN_7; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_185 = 3'h1 == head ? io_decoder_0_entry_sourceTag2_threadId : _GEN_67; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_186 = 3'h2 == head ? io_decoder_0_entry_sourceTag2_threadId : _GEN_22; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_187 = 3'h3 == head ? io_decoder_0_entry_sourceTag2_threadId : _GEN_82; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_188 = 3'h4 == head ? io_decoder_0_entry_sourceTag2_threadId : _GEN_37; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_189 = 3'h5 == head ? io_decoder_0_entry_sourceTag2_threadId : _GEN_97; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_190 = 3'h6 == head ? io_decoder_0_entry_sourceTag2_threadId : _GEN_52; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_191 = 3'h7 == head ? io_decoder_0_entry_sourceTag2_threadId : _GEN_112; // @[ReservationStation.scala 69:{31,31}]
  wire [3:0] _GEN_192 = 3'h0 == head ? io_decoder_0_entry_sourceTag2_id : _GEN_6; // @[ReservationStation.scala 69:{31,31}]
  wire [3:0] _GEN_193 = 3'h1 == head ? io_decoder_0_entry_sourceTag2_id : _GEN_66; // @[ReservationStation.scala 69:{31,31}]
  wire [3:0] _GEN_194 = 3'h2 == head ? io_decoder_0_entry_sourceTag2_id : _GEN_21; // @[ReservationStation.scala 69:{31,31}]
  wire [3:0] _GEN_195 = 3'h3 == head ? io_decoder_0_entry_sourceTag2_id : _GEN_81; // @[ReservationStation.scala 69:{31,31}]
  wire [3:0] _GEN_196 = 3'h4 == head ? io_decoder_0_entry_sourceTag2_id : _GEN_36; // @[ReservationStation.scala 69:{31,31}]
  wire [3:0] _GEN_197 = 3'h5 == head ? io_decoder_0_entry_sourceTag2_id : _GEN_96; // @[ReservationStation.scala 69:{31,31}]
  wire [3:0] _GEN_198 = 3'h6 == head ? io_decoder_0_entry_sourceTag2_id : _GEN_51; // @[ReservationStation.scala 69:{31,31}]
  wire [3:0] _GEN_199 = 3'h7 == head ? io_decoder_0_entry_sourceTag2_id : _GEN_111; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_200 = 3'h0 == head ? io_decoder_0_entry_ready2 : _GEN_5; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_201 = 3'h1 == head ? io_decoder_0_entry_ready2 : _GEN_65; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_202 = 3'h2 == head ? io_decoder_0_entry_ready2 : _GEN_20; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_203 = 3'h3 == head ? io_decoder_0_entry_ready2 : _GEN_80; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_204 = 3'h4 == head ? io_decoder_0_entry_ready2 : _GEN_35; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_205 = 3'h5 == head ? io_decoder_0_entry_ready2 : _GEN_95; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_206 = 3'h6 == head ? io_decoder_0_entry_ready2 : _GEN_50; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_207 = 3'h7 == head ? io_decoder_0_entry_ready2 : _GEN_110; // @[ReservationStation.scala 69:{31,31}]
  wire [63:0] _GEN_208 = 3'h0 == head ? io_decoder_0_entry_value2 : _GEN_4; // @[ReservationStation.scala 69:{31,31}]
  wire [63:0] _GEN_209 = 3'h1 == head ? io_decoder_0_entry_value2 : _GEN_64; // @[ReservationStation.scala 69:{31,31}]
  wire [63:0] _GEN_210 = 3'h2 == head ? io_decoder_0_entry_value2 : _GEN_19; // @[ReservationStation.scala 69:{31,31}]
  wire [63:0] _GEN_211 = 3'h3 == head ? io_decoder_0_entry_value2 : _GEN_79; // @[ReservationStation.scala 69:{31,31}]
  wire [63:0] _GEN_212 = 3'h4 == head ? io_decoder_0_entry_value2 : _GEN_34; // @[ReservationStation.scala 69:{31,31}]
  wire [63:0] _GEN_213 = 3'h5 == head ? io_decoder_0_entry_value2 : _GEN_94; // @[ReservationStation.scala 69:{31,31}]
  wire [63:0] _GEN_214 = 3'h6 == head ? io_decoder_0_entry_value2 : _GEN_49; // @[ReservationStation.scala 69:{31,31}]
  wire [63:0] _GEN_215 = 3'h7 == head ? io_decoder_0_entry_value2 : _GEN_109; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_216 = 3'h0 == head ? 1'h0 : _GEN_3; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_217 = 3'h1 == head ? 1'h0 : _GEN_63; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_218 = 3'h2 == head ? 1'h0 : _GEN_18; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_219 = 3'h3 == head ? 1'h0 : _GEN_78; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_220 = 3'h4 == head ? 1'h0 : _GEN_33; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_221 = 3'h5 == head ? 1'h0 : _GEN_93; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_222 = 3'h6 == head ? 1'h0 : _GEN_48; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_223 = 3'h7 == head ? 1'h0 : _GEN_108; // @[ReservationStation.scala 69:{31,31}]
  wire [3:0] _GEN_224 = 3'h0 == head ? io_decoder_0_entry_destinationTag_id : _GEN_2; // @[ReservationStation.scala 69:{31,31}]
  wire [3:0] _GEN_225 = 3'h1 == head ? io_decoder_0_entry_destinationTag_id : _GEN_62; // @[ReservationStation.scala 69:{31,31}]
  wire [3:0] _GEN_226 = 3'h2 == head ? io_decoder_0_entry_destinationTag_id : _GEN_17; // @[ReservationStation.scala 69:{31,31}]
  wire [3:0] _GEN_227 = 3'h3 == head ? io_decoder_0_entry_destinationTag_id : _GEN_77; // @[ReservationStation.scala 69:{31,31}]
  wire [3:0] _GEN_228 = 3'h4 == head ? io_decoder_0_entry_destinationTag_id : _GEN_32; // @[ReservationStation.scala 69:{31,31}]
  wire [3:0] _GEN_229 = 3'h5 == head ? io_decoder_0_entry_destinationTag_id : _GEN_92; // @[ReservationStation.scala 69:{31,31}]
  wire [3:0] _GEN_230 = 3'h6 == head ? io_decoder_0_entry_destinationTag_id : _GEN_47; // @[ReservationStation.scala 69:{31,31}]
  wire [3:0] _GEN_231 = 3'h7 == head ? io_decoder_0_entry_destinationTag_id : _GEN_107; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_232 = 3'h0 == head ? io_decoder_0_entry_wasCompressed : _GEN_1; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_233 = 3'h1 == head ? io_decoder_0_entry_wasCompressed : _GEN_61; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_234 = 3'h2 == head ? io_decoder_0_entry_wasCompressed : _GEN_16; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_235 = 3'h3 == head ? io_decoder_0_entry_wasCompressed : _GEN_76; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_236 = 3'h4 == head ? io_decoder_0_entry_wasCompressed : _GEN_31; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_237 = 3'h5 == head ? io_decoder_0_entry_wasCompressed : _GEN_91; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_238 = 3'h6 == head ? io_decoder_0_entry_wasCompressed : _GEN_46; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_239 = 3'h7 == head ? io_decoder_0_entry_wasCompressed : _GEN_106; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_240 = 3'h0 == head ? io_decoder_0_entry_valid : _GEN_0; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_241 = 3'h1 == head ? io_decoder_0_entry_valid : _GEN_60; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_242 = 3'h2 == head ? io_decoder_0_entry_valid : _GEN_15; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_243 = 3'h3 == head ? io_decoder_0_entry_valid : _GEN_75; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_244 = 3'h4 == head ? io_decoder_0_entry_valid : _GEN_30; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_245 = 3'h5 == head ? io_decoder_0_entry_valid : _GEN_90; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_246 = 3'h6 == head ? io_decoder_0_entry_valid : _GEN_45; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_247 = 3'h7 == head ? io_decoder_0_entry_valid : _GEN_105; // @[ReservationStation.scala 69:{31,31}]
  wire [6:0] _GEN_248 = io_decoder_0_entry_valid ? _GEN_128 : _GEN_14; // @[ReservationStation.scala 68:39]
  wire [6:0] _GEN_249 = io_decoder_0_entry_valid ? _GEN_129 : _GEN_74; // @[ReservationStation.scala 68:39]
  wire [6:0] _GEN_250 = io_decoder_0_entry_valid ? _GEN_130 : _GEN_29; // @[ReservationStation.scala 68:39]
  wire [6:0] _GEN_251 = io_decoder_0_entry_valid ? _GEN_131 : _GEN_89; // @[ReservationStation.scala 68:39]
  wire [6:0] _GEN_252 = io_decoder_0_entry_valid ? _GEN_132 : _GEN_44; // @[ReservationStation.scala 68:39]
  wire [6:0] _GEN_253 = io_decoder_0_entry_valid ? _GEN_133 : _GEN_104; // @[ReservationStation.scala 68:39]
  wire [6:0] _GEN_254 = io_decoder_0_entry_valid ? _GEN_134 : _GEN_59; // @[ReservationStation.scala 68:39]
  wire [6:0] _GEN_255 = io_decoder_0_entry_valid ? _GEN_135 : _GEN_119; // @[ReservationStation.scala 68:39]
  wire [2:0] _GEN_256 = io_decoder_0_entry_valid ? _GEN_136 : _GEN_13; // @[ReservationStation.scala 68:39]
  wire [2:0] _GEN_257 = io_decoder_0_entry_valid ? _GEN_137 : _GEN_73; // @[ReservationStation.scala 68:39]
  wire [2:0] _GEN_258 = io_decoder_0_entry_valid ? _GEN_138 : _GEN_28; // @[ReservationStation.scala 68:39]
  wire [2:0] _GEN_259 = io_decoder_0_entry_valid ? _GEN_139 : _GEN_88; // @[ReservationStation.scala 68:39]
  wire [2:0] _GEN_260 = io_decoder_0_entry_valid ? _GEN_140 : _GEN_43; // @[ReservationStation.scala 68:39]
  wire [2:0] _GEN_261 = io_decoder_0_entry_valid ? _GEN_141 : _GEN_103; // @[ReservationStation.scala 68:39]
  wire [2:0] _GEN_262 = io_decoder_0_entry_valid ? _GEN_142 : _GEN_58; // @[ReservationStation.scala 68:39]
  wire [2:0] _GEN_263 = io_decoder_0_entry_valid ? _GEN_143 : _GEN_118; // @[ReservationStation.scala 68:39]
  wire [11:0] _GEN_264 = io_decoder_0_entry_valid ? _GEN_144 : _GEN_12; // @[ReservationStation.scala 68:39]
  wire [11:0] _GEN_265 = io_decoder_0_entry_valid ? _GEN_145 : _GEN_72; // @[ReservationStation.scala 68:39]
  wire [11:0] _GEN_266 = io_decoder_0_entry_valid ? _GEN_146 : _GEN_27; // @[ReservationStation.scala 68:39]
  wire [11:0] _GEN_267 = io_decoder_0_entry_valid ? _GEN_147 : _GEN_87; // @[ReservationStation.scala 68:39]
  wire [11:0] _GEN_268 = io_decoder_0_entry_valid ? _GEN_148 : _GEN_42; // @[ReservationStation.scala 68:39]
  wire [11:0] _GEN_269 = io_decoder_0_entry_valid ? _GEN_149 : _GEN_102; // @[ReservationStation.scala 68:39]
  wire [11:0] _GEN_270 = io_decoder_0_entry_valid ? _GEN_150 : _GEN_57; // @[ReservationStation.scala 68:39]
  wire [11:0] _GEN_271 = io_decoder_0_entry_valid ? _GEN_151 : _GEN_117; // @[ReservationStation.scala 68:39]
  wire  _GEN_272 = io_decoder_0_entry_valid ? _GEN_152 : _GEN_11; // @[ReservationStation.scala 68:39]
  wire  _GEN_273 = io_decoder_0_entry_valid ? _GEN_153 : _GEN_71; // @[ReservationStation.scala 68:39]
  wire  _GEN_274 = io_decoder_0_entry_valid ? _GEN_154 : _GEN_26; // @[ReservationStation.scala 68:39]
  wire  _GEN_275 = io_decoder_0_entry_valid ? _GEN_155 : _GEN_86; // @[ReservationStation.scala 68:39]
  wire  _GEN_276 = io_decoder_0_entry_valid ? _GEN_156 : _GEN_41; // @[ReservationStation.scala 68:39]
  wire  _GEN_277 = io_decoder_0_entry_valid ? _GEN_157 : _GEN_101; // @[ReservationStation.scala 68:39]
  wire  _GEN_278 = io_decoder_0_entry_valid ? _GEN_158 : _GEN_56; // @[ReservationStation.scala 68:39]
  wire  _GEN_279 = io_decoder_0_entry_valid ? _GEN_159 : _GEN_116; // @[ReservationStation.scala 68:39]
  wire [3:0] _GEN_280 = io_decoder_0_entry_valid ? _GEN_160 : _GEN_10; // @[ReservationStation.scala 68:39]
  wire [3:0] _GEN_281 = io_decoder_0_entry_valid ? _GEN_161 : _GEN_70; // @[ReservationStation.scala 68:39]
  wire [3:0] _GEN_282 = io_decoder_0_entry_valid ? _GEN_162 : _GEN_25; // @[ReservationStation.scala 68:39]
  wire [3:0] _GEN_283 = io_decoder_0_entry_valid ? _GEN_163 : _GEN_85; // @[ReservationStation.scala 68:39]
  wire [3:0] _GEN_284 = io_decoder_0_entry_valid ? _GEN_164 : _GEN_40; // @[ReservationStation.scala 68:39]
  wire [3:0] _GEN_285 = io_decoder_0_entry_valid ? _GEN_165 : _GEN_100; // @[ReservationStation.scala 68:39]
  wire [3:0] _GEN_286 = io_decoder_0_entry_valid ? _GEN_166 : _GEN_55; // @[ReservationStation.scala 68:39]
  wire [3:0] _GEN_287 = io_decoder_0_entry_valid ? _GEN_167 : _GEN_115; // @[ReservationStation.scala 68:39]
  wire  _GEN_288 = io_decoder_0_entry_valid ? _GEN_168 : _GEN_9; // @[ReservationStation.scala 68:39]
  wire  _GEN_289 = io_decoder_0_entry_valid ? _GEN_169 : _GEN_69; // @[ReservationStation.scala 68:39]
  wire  _GEN_290 = io_decoder_0_entry_valid ? _GEN_170 : _GEN_24; // @[ReservationStation.scala 68:39]
  wire  _GEN_291 = io_decoder_0_entry_valid ? _GEN_171 : _GEN_84; // @[ReservationStation.scala 68:39]
  wire  _GEN_292 = io_decoder_0_entry_valid ? _GEN_172 : _GEN_39; // @[ReservationStation.scala 68:39]
  wire  _GEN_293 = io_decoder_0_entry_valid ? _GEN_173 : _GEN_99; // @[ReservationStation.scala 68:39]
  wire  _GEN_294 = io_decoder_0_entry_valid ? _GEN_174 : _GEN_54; // @[ReservationStation.scala 68:39]
  wire  _GEN_295 = io_decoder_0_entry_valid ? _GEN_175 : _GEN_114; // @[ReservationStation.scala 68:39]
  wire [63:0] _GEN_296 = io_decoder_0_entry_valid ? _GEN_176 : _GEN_8; // @[ReservationStation.scala 68:39]
  wire [63:0] _GEN_297 = io_decoder_0_entry_valid ? _GEN_177 : _GEN_68; // @[ReservationStation.scala 68:39]
  wire [63:0] _GEN_298 = io_decoder_0_entry_valid ? _GEN_178 : _GEN_23; // @[ReservationStation.scala 68:39]
  wire [63:0] _GEN_299 = io_decoder_0_entry_valid ? _GEN_179 : _GEN_83; // @[ReservationStation.scala 68:39]
  wire [63:0] _GEN_300 = io_decoder_0_entry_valid ? _GEN_180 : _GEN_38; // @[ReservationStation.scala 68:39]
  wire [63:0] _GEN_301 = io_decoder_0_entry_valid ? _GEN_181 : _GEN_98; // @[ReservationStation.scala 68:39]
  wire [63:0] _GEN_302 = io_decoder_0_entry_valid ? _GEN_182 : _GEN_53; // @[ReservationStation.scala 68:39]
  wire [63:0] _GEN_303 = io_decoder_0_entry_valid ? _GEN_183 : _GEN_113; // @[ReservationStation.scala 68:39]
  wire  _GEN_304 = io_decoder_0_entry_valid ? _GEN_184 : _GEN_7; // @[ReservationStation.scala 68:39]
  wire  _GEN_305 = io_decoder_0_entry_valid ? _GEN_185 : _GEN_67; // @[ReservationStation.scala 68:39]
  wire  _GEN_306 = io_decoder_0_entry_valid ? _GEN_186 : _GEN_22; // @[ReservationStation.scala 68:39]
  wire  _GEN_307 = io_decoder_0_entry_valid ? _GEN_187 : _GEN_82; // @[ReservationStation.scala 68:39]
  wire  _GEN_308 = io_decoder_0_entry_valid ? _GEN_188 : _GEN_37; // @[ReservationStation.scala 68:39]
  wire  _GEN_309 = io_decoder_0_entry_valid ? _GEN_189 : _GEN_97; // @[ReservationStation.scala 68:39]
  wire  _GEN_310 = io_decoder_0_entry_valid ? _GEN_190 : _GEN_52; // @[ReservationStation.scala 68:39]
  wire  _GEN_311 = io_decoder_0_entry_valid ? _GEN_191 : _GEN_112; // @[ReservationStation.scala 68:39]
  wire [3:0] _GEN_312 = io_decoder_0_entry_valid ? _GEN_192 : _GEN_6; // @[ReservationStation.scala 68:39]
  wire [3:0] _GEN_313 = io_decoder_0_entry_valid ? _GEN_193 : _GEN_66; // @[ReservationStation.scala 68:39]
  wire [3:0] _GEN_314 = io_decoder_0_entry_valid ? _GEN_194 : _GEN_21; // @[ReservationStation.scala 68:39]
  wire [3:0] _GEN_315 = io_decoder_0_entry_valid ? _GEN_195 : _GEN_81; // @[ReservationStation.scala 68:39]
  wire [3:0] _GEN_316 = io_decoder_0_entry_valid ? _GEN_196 : _GEN_36; // @[ReservationStation.scala 68:39]
  wire [3:0] _GEN_317 = io_decoder_0_entry_valid ? _GEN_197 : _GEN_96; // @[ReservationStation.scala 68:39]
  wire [3:0] _GEN_318 = io_decoder_0_entry_valid ? _GEN_198 : _GEN_51; // @[ReservationStation.scala 68:39]
  wire [3:0] _GEN_319 = io_decoder_0_entry_valid ? _GEN_199 : _GEN_111; // @[ReservationStation.scala 68:39]
  wire  _GEN_320 = io_decoder_0_entry_valid ? _GEN_200 : _GEN_5; // @[ReservationStation.scala 68:39]
  wire  _GEN_321 = io_decoder_0_entry_valid ? _GEN_201 : _GEN_65; // @[ReservationStation.scala 68:39]
  wire  _GEN_322 = io_decoder_0_entry_valid ? _GEN_202 : _GEN_20; // @[ReservationStation.scala 68:39]
  wire  _GEN_323 = io_decoder_0_entry_valid ? _GEN_203 : _GEN_80; // @[ReservationStation.scala 68:39]
  wire  _GEN_324 = io_decoder_0_entry_valid ? _GEN_204 : _GEN_35; // @[ReservationStation.scala 68:39]
  wire  _GEN_325 = io_decoder_0_entry_valid ? _GEN_205 : _GEN_95; // @[ReservationStation.scala 68:39]
  wire  _GEN_326 = io_decoder_0_entry_valid ? _GEN_206 : _GEN_50; // @[ReservationStation.scala 68:39]
  wire  _GEN_327 = io_decoder_0_entry_valid ? _GEN_207 : _GEN_110; // @[ReservationStation.scala 68:39]
  wire [63:0] _GEN_328 = io_decoder_0_entry_valid ? _GEN_208 : _GEN_4; // @[ReservationStation.scala 68:39]
  wire [63:0] _GEN_329 = io_decoder_0_entry_valid ? _GEN_209 : _GEN_64; // @[ReservationStation.scala 68:39]
  wire [63:0] _GEN_330 = io_decoder_0_entry_valid ? _GEN_210 : _GEN_19; // @[ReservationStation.scala 68:39]
  wire [63:0] _GEN_331 = io_decoder_0_entry_valid ? _GEN_211 : _GEN_79; // @[ReservationStation.scala 68:39]
  wire [63:0] _GEN_332 = io_decoder_0_entry_valid ? _GEN_212 : _GEN_34; // @[ReservationStation.scala 68:39]
  wire [63:0] _GEN_333 = io_decoder_0_entry_valid ? _GEN_213 : _GEN_94; // @[ReservationStation.scala 68:39]
  wire [63:0] _GEN_334 = io_decoder_0_entry_valid ? _GEN_214 : _GEN_49; // @[ReservationStation.scala 68:39]
  wire [63:0] _GEN_335 = io_decoder_0_entry_valid ? _GEN_215 : _GEN_109; // @[ReservationStation.scala 68:39]
  wire  _GEN_336 = io_decoder_0_entry_valid ? _GEN_216 : _GEN_3; // @[ReservationStation.scala 68:39]
  wire  _GEN_337 = io_decoder_0_entry_valid ? _GEN_217 : _GEN_63; // @[ReservationStation.scala 68:39]
  wire  _GEN_338 = io_decoder_0_entry_valid ? _GEN_218 : _GEN_18; // @[ReservationStation.scala 68:39]
  wire  _GEN_339 = io_decoder_0_entry_valid ? _GEN_219 : _GEN_78; // @[ReservationStation.scala 68:39]
  wire  _GEN_340 = io_decoder_0_entry_valid ? _GEN_220 : _GEN_33; // @[ReservationStation.scala 68:39]
  wire  _GEN_341 = io_decoder_0_entry_valid ? _GEN_221 : _GEN_93; // @[ReservationStation.scala 68:39]
  wire  _GEN_342 = io_decoder_0_entry_valid ? _GEN_222 : _GEN_48; // @[ReservationStation.scala 68:39]
  wire  _GEN_343 = io_decoder_0_entry_valid ? _GEN_223 : _GEN_108; // @[ReservationStation.scala 68:39]
  wire [3:0] _GEN_344 = io_decoder_0_entry_valid ? _GEN_224 : _GEN_2; // @[ReservationStation.scala 68:39]
  wire [3:0] _GEN_345 = io_decoder_0_entry_valid ? _GEN_225 : _GEN_62; // @[ReservationStation.scala 68:39]
  wire [3:0] _GEN_346 = io_decoder_0_entry_valid ? _GEN_226 : _GEN_17; // @[ReservationStation.scala 68:39]
  wire [3:0] _GEN_347 = io_decoder_0_entry_valid ? _GEN_227 : _GEN_77; // @[ReservationStation.scala 68:39]
  wire [3:0] _GEN_348 = io_decoder_0_entry_valid ? _GEN_228 : _GEN_32; // @[ReservationStation.scala 68:39]
  wire [3:0] _GEN_349 = io_decoder_0_entry_valid ? _GEN_229 : _GEN_92; // @[ReservationStation.scala 68:39]
  wire [3:0] _GEN_350 = io_decoder_0_entry_valid ? _GEN_230 : _GEN_47; // @[ReservationStation.scala 68:39]
  wire [3:0] _GEN_351 = io_decoder_0_entry_valid ? _GEN_231 : _GEN_107; // @[ReservationStation.scala 68:39]
  wire  _GEN_352 = io_decoder_0_entry_valid ? _GEN_232 : _GEN_1; // @[ReservationStation.scala 68:39]
  wire  _GEN_353 = io_decoder_0_entry_valid ? _GEN_233 : _GEN_61; // @[ReservationStation.scala 68:39]
  wire  _GEN_354 = io_decoder_0_entry_valid ? _GEN_234 : _GEN_16; // @[ReservationStation.scala 68:39]
  wire  _GEN_355 = io_decoder_0_entry_valid ? _GEN_235 : _GEN_76; // @[ReservationStation.scala 68:39]
  wire  _GEN_356 = io_decoder_0_entry_valid ? _GEN_236 : _GEN_31; // @[ReservationStation.scala 68:39]
  wire  _GEN_357 = io_decoder_0_entry_valid ? _GEN_237 : _GEN_91; // @[ReservationStation.scala 68:39]
  wire  _GEN_358 = io_decoder_0_entry_valid ? _GEN_238 : _GEN_46; // @[ReservationStation.scala 68:39]
  wire  _GEN_359 = io_decoder_0_entry_valid ? _GEN_239 : _GEN_106; // @[ReservationStation.scala 68:39]
  wire  _GEN_360 = io_decoder_0_entry_valid ? _GEN_240 : _GEN_0; // @[ReservationStation.scala 68:39]
  wire  _GEN_361 = io_decoder_0_entry_valid ? _GEN_241 : _GEN_60; // @[ReservationStation.scala 68:39]
  wire  _GEN_362 = io_decoder_0_entry_valid ? _GEN_242 : _GEN_15; // @[ReservationStation.scala 68:39]
  wire  _GEN_363 = io_decoder_0_entry_valid ? _GEN_243 : _GEN_75; // @[ReservationStation.scala 68:39]
  wire  _GEN_364 = io_decoder_0_entry_valid ? _GEN_244 : _GEN_30; // @[ReservationStation.scala 68:39]
  wire  _GEN_365 = io_decoder_0_entry_valid ? _GEN_245 : _GEN_90; // @[ReservationStation.scala 68:39]
  wire  _GEN_366 = io_decoder_0_entry_valid ? _GEN_246 : _GEN_45; // @[ReservationStation.scala 68:39]
  wire  _GEN_367 = io_decoder_0_entry_valid ? _GEN_247 : _GEN_105; // @[ReservationStation.scala 68:39]
  wire [6:0] _GEN_369 = ~_GEN_127 ? _GEN_248 : _GEN_14; // @[ReservationStation.scala 66:40]
  wire [6:0] _GEN_370 = ~_GEN_127 ? _GEN_249 : _GEN_74; // @[ReservationStation.scala 66:40]
  wire [6:0] _GEN_371 = ~_GEN_127 ? _GEN_250 : _GEN_29; // @[ReservationStation.scala 66:40]
  wire [6:0] _GEN_372 = ~_GEN_127 ? _GEN_251 : _GEN_89; // @[ReservationStation.scala 66:40]
  wire [6:0] _GEN_373 = ~_GEN_127 ? _GEN_252 : _GEN_44; // @[ReservationStation.scala 66:40]
  wire [6:0] _GEN_374 = ~_GEN_127 ? _GEN_253 : _GEN_104; // @[ReservationStation.scala 66:40]
  wire [6:0] _GEN_375 = ~_GEN_127 ? _GEN_254 : _GEN_59; // @[ReservationStation.scala 66:40]
  wire [6:0] _GEN_376 = ~_GEN_127 ? _GEN_255 : _GEN_119; // @[ReservationStation.scala 66:40]
  wire [2:0] _GEN_377 = ~_GEN_127 ? _GEN_256 : _GEN_13; // @[ReservationStation.scala 66:40]
  wire [2:0] _GEN_378 = ~_GEN_127 ? _GEN_257 : _GEN_73; // @[ReservationStation.scala 66:40]
  wire [2:0] _GEN_379 = ~_GEN_127 ? _GEN_258 : _GEN_28; // @[ReservationStation.scala 66:40]
  wire [2:0] _GEN_380 = ~_GEN_127 ? _GEN_259 : _GEN_88; // @[ReservationStation.scala 66:40]
  wire [2:0] _GEN_381 = ~_GEN_127 ? _GEN_260 : _GEN_43; // @[ReservationStation.scala 66:40]
  wire [2:0] _GEN_382 = ~_GEN_127 ? _GEN_261 : _GEN_103; // @[ReservationStation.scala 66:40]
  wire [2:0] _GEN_383 = ~_GEN_127 ? _GEN_262 : _GEN_58; // @[ReservationStation.scala 66:40]
  wire [2:0] _GEN_384 = ~_GEN_127 ? _GEN_263 : _GEN_118; // @[ReservationStation.scala 66:40]
  wire [11:0] _GEN_385 = ~_GEN_127 ? _GEN_264 : _GEN_12; // @[ReservationStation.scala 66:40]
  wire [11:0] _GEN_386 = ~_GEN_127 ? _GEN_265 : _GEN_72; // @[ReservationStation.scala 66:40]
  wire [11:0] _GEN_387 = ~_GEN_127 ? _GEN_266 : _GEN_27; // @[ReservationStation.scala 66:40]
  wire [11:0] _GEN_388 = ~_GEN_127 ? _GEN_267 : _GEN_87; // @[ReservationStation.scala 66:40]
  wire [11:0] _GEN_389 = ~_GEN_127 ? _GEN_268 : _GEN_42; // @[ReservationStation.scala 66:40]
  wire [11:0] _GEN_390 = ~_GEN_127 ? _GEN_269 : _GEN_102; // @[ReservationStation.scala 66:40]
  wire [11:0] _GEN_391 = ~_GEN_127 ? _GEN_270 : _GEN_57; // @[ReservationStation.scala 66:40]
  wire [11:0] _GEN_392 = ~_GEN_127 ? _GEN_271 : _GEN_117; // @[ReservationStation.scala 66:40]
  wire  _GEN_393 = ~_GEN_127 ? _GEN_272 : _GEN_11; // @[ReservationStation.scala 66:40]
  wire  _GEN_394 = ~_GEN_127 ? _GEN_273 : _GEN_71; // @[ReservationStation.scala 66:40]
  wire  _GEN_395 = ~_GEN_127 ? _GEN_274 : _GEN_26; // @[ReservationStation.scala 66:40]
  wire  _GEN_396 = ~_GEN_127 ? _GEN_275 : _GEN_86; // @[ReservationStation.scala 66:40]
  wire  _GEN_397 = ~_GEN_127 ? _GEN_276 : _GEN_41; // @[ReservationStation.scala 66:40]
  wire  _GEN_398 = ~_GEN_127 ? _GEN_277 : _GEN_101; // @[ReservationStation.scala 66:40]
  wire  _GEN_399 = ~_GEN_127 ? _GEN_278 : _GEN_56; // @[ReservationStation.scala 66:40]
  wire  _GEN_400 = ~_GEN_127 ? _GEN_279 : _GEN_116; // @[ReservationStation.scala 66:40]
  wire [3:0] _GEN_401 = ~_GEN_127 ? _GEN_280 : _GEN_10; // @[ReservationStation.scala 66:40]
  wire [3:0] _GEN_402 = ~_GEN_127 ? _GEN_281 : _GEN_70; // @[ReservationStation.scala 66:40]
  wire [3:0] _GEN_403 = ~_GEN_127 ? _GEN_282 : _GEN_25; // @[ReservationStation.scala 66:40]
  wire [3:0] _GEN_404 = ~_GEN_127 ? _GEN_283 : _GEN_85; // @[ReservationStation.scala 66:40]
  wire [3:0] _GEN_405 = ~_GEN_127 ? _GEN_284 : _GEN_40; // @[ReservationStation.scala 66:40]
  wire [3:0] _GEN_406 = ~_GEN_127 ? _GEN_285 : _GEN_100; // @[ReservationStation.scala 66:40]
  wire [3:0] _GEN_407 = ~_GEN_127 ? _GEN_286 : _GEN_55; // @[ReservationStation.scala 66:40]
  wire [3:0] _GEN_408 = ~_GEN_127 ? _GEN_287 : _GEN_115; // @[ReservationStation.scala 66:40]
  wire  _GEN_409 = ~_GEN_127 ? _GEN_288 : _GEN_9; // @[ReservationStation.scala 66:40]
  wire  _GEN_410 = ~_GEN_127 ? _GEN_289 : _GEN_69; // @[ReservationStation.scala 66:40]
  wire  _GEN_411 = ~_GEN_127 ? _GEN_290 : _GEN_24; // @[ReservationStation.scala 66:40]
  wire  _GEN_412 = ~_GEN_127 ? _GEN_291 : _GEN_84; // @[ReservationStation.scala 66:40]
  wire  _GEN_413 = ~_GEN_127 ? _GEN_292 : _GEN_39; // @[ReservationStation.scala 66:40]
  wire  _GEN_414 = ~_GEN_127 ? _GEN_293 : _GEN_99; // @[ReservationStation.scala 66:40]
  wire  _GEN_415 = ~_GEN_127 ? _GEN_294 : _GEN_54; // @[ReservationStation.scala 66:40]
  wire  _GEN_416 = ~_GEN_127 ? _GEN_295 : _GEN_114; // @[ReservationStation.scala 66:40]
  wire [63:0] _GEN_417 = ~_GEN_127 ? _GEN_296 : _GEN_8; // @[ReservationStation.scala 66:40]
  wire [63:0] _GEN_418 = ~_GEN_127 ? _GEN_297 : _GEN_68; // @[ReservationStation.scala 66:40]
  wire [63:0] _GEN_419 = ~_GEN_127 ? _GEN_298 : _GEN_23; // @[ReservationStation.scala 66:40]
  wire [63:0] _GEN_420 = ~_GEN_127 ? _GEN_299 : _GEN_83; // @[ReservationStation.scala 66:40]
  wire [63:0] _GEN_421 = ~_GEN_127 ? _GEN_300 : _GEN_38; // @[ReservationStation.scala 66:40]
  wire [63:0] _GEN_422 = ~_GEN_127 ? _GEN_301 : _GEN_98; // @[ReservationStation.scala 66:40]
  wire [63:0] _GEN_423 = ~_GEN_127 ? _GEN_302 : _GEN_53; // @[ReservationStation.scala 66:40]
  wire [63:0] _GEN_424 = ~_GEN_127 ? _GEN_303 : _GEN_113; // @[ReservationStation.scala 66:40]
  wire  _GEN_425 = ~_GEN_127 ? _GEN_304 : _GEN_7; // @[ReservationStation.scala 66:40]
  wire  _GEN_426 = ~_GEN_127 ? _GEN_305 : _GEN_67; // @[ReservationStation.scala 66:40]
  wire  _GEN_427 = ~_GEN_127 ? _GEN_306 : _GEN_22; // @[ReservationStation.scala 66:40]
  wire  _GEN_428 = ~_GEN_127 ? _GEN_307 : _GEN_82; // @[ReservationStation.scala 66:40]
  wire  _GEN_429 = ~_GEN_127 ? _GEN_308 : _GEN_37; // @[ReservationStation.scala 66:40]
  wire  _GEN_430 = ~_GEN_127 ? _GEN_309 : _GEN_97; // @[ReservationStation.scala 66:40]
  wire  _GEN_431 = ~_GEN_127 ? _GEN_310 : _GEN_52; // @[ReservationStation.scala 66:40]
  wire  _GEN_432 = ~_GEN_127 ? _GEN_311 : _GEN_112; // @[ReservationStation.scala 66:40]
  wire [3:0] _GEN_433 = ~_GEN_127 ? _GEN_312 : _GEN_6; // @[ReservationStation.scala 66:40]
  wire [3:0] _GEN_434 = ~_GEN_127 ? _GEN_313 : _GEN_66; // @[ReservationStation.scala 66:40]
  wire [3:0] _GEN_435 = ~_GEN_127 ? _GEN_314 : _GEN_21; // @[ReservationStation.scala 66:40]
  wire [3:0] _GEN_436 = ~_GEN_127 ? _GEN_315 : _GEN_81; // @[ReservationStation.scala 66:40]
  wire [3:0] _GEN_437 = ~_GEN_127 ? _GEN_316 : _GEN_36; // @[ReservationStation.scala 66:40]
  wire [3:0] _GEN_438 = ~_GEN_127 ? _GEN_317 : _GEN_96; // @[ReservationStation.scala 66:40]
  wire [3:0] _GEN_439 = ~_GEN_127 ? _GEN_318 : _GEN_51; // @[ReservationStation.scala 66:40]
  wire [3:0] _GEN_440 = ~_GEN_127 ? _GEN_319 : _GEN_111; // @[ReservationStation.scala 66:40]
  wire  _GEN_441 = ~_GEN_127 ? _GEN_320 : _GEN_5; // @[ReservationStation.scala 66:40]
  wire  _GEN_442 = ~_GEN_127 ? _GEN_321 : _GEN_65; // @[ReservationStation.scala 66:40]
  wire  _GEN_443 = ~_GEN_127 ? _GEN_322 : _GEN_20; // @[ReservationStation.scala 66:40]
  wire  _GEN_444 = ~_GEN_127 ? _GEN_323 : _GEN_80; // @[ReservationStation.scala 66:40]
  wire  _GEN_445 = ~_GEN_127 ? _GEN_324 : _GEN_35; // @[ReservationStation.scala 66:40]
  wire  _GEN_446 = ~_GEN_127 ? _GEN_325 : _GEN_95; // @[ReservationStation.scala 66:40]
  wire  _GEN_447 = ~_GEN_127 ? _GEN_326 : _GEN_50; // @[ReservationStation.scala 66:40]
  wire  _GEN_448 = ~_GEN_127 ? _GEN_327 : _GEN_110; // @[ReservationStation.scala 66:40]
  wire [63:0] _GEN_449 = ~_GEN_127 ? _GEN_328 : _GEN_4; // @[ReservationStation.scala 66:40]
  wire [63:0] _GEN_450 = ~_GEN_127 ? _GEN_329 : _GEN_64; // @[ReservationStation.scala 66:40]
  wire [63:0] _GEN_451 = ~_GEN_127 ? _GEN_330 : _GEN_19; // @[ReservationStation.scala 66:40]
  wire [63:0] _GEN_452 = ~_GEN_127 ? _GEN_331 : _GEN_79; // @[ReservationStation.scala 66:40]
  wire [63:0] _GEN_453 = ~_GEN_127 ? _GEN_332 : _GEN_34; // @[ReservationStation.scala 66:40]
  wire [63:0] _GEN_454 = ~_GEN_127 ? _GEN_333 : _GEN_94; // @[ReservationStation.scala 66:40]
  wire [63:0] _GEN_455 = ~_GEN_127 ? _GEN_334 : _GEN_49; // @[ReservationStation.scala 66:40]
  wire [63:0] _GEN_456 = ~_GEN_127 ? _GEN_335 : _GEN_109; // @[ReservationStation.scala 66:40]
  wire  _GEN_457 = ~_GEN_127 ? _GEN_336 : _GEN_3; // @[ReservationStation.scala 66:40]
  wire  _GEN_458 = ~_GEN_127 ? _GEN_337 : _GEN_63; // @[ReservationStation.scala 66:40]
  wire  _GEN_459 = ~_GEN_127 ? _GEN_338 : _GEN_18; // @[ReservationStation.scala 66:40]
  wire  _GEN_460 = ~_GEN_127 ? _GEN_339 : _GEN_78; // @[ReservationStation.scala 66:40]
  wire  _GEN_461 = ~_GEN_127 ? _GEN_340 : _GEN_33; // @[ReservationStation.scala 66:40]
  wire  _GEN_462 = ~_GEN_127 ? _GEN_341 : _GEN_93; // @[ReservationStation.scala 66:40]
  wire  _GEN_463 = ~_GEN_127 ? _GEN_342 : _GEN_48; // @[ReservationStation.scala 66:40]
  wire  _GEN_464 = ~_GEN_127 ? _GEN_343 : _GEN_108; // @[ReservationStation.scala 66:40]
  wire [3:0] _GEN_465 = ~_GEN_127 ? _GEN_344 : _GEN_2; // @[ReservationStation.scala 66:40]
  wire [3:0] _GEN_466 = ~_GEN_127 ? _GEN_345 : _GEN_62; // @[ReservationStation.scala 66:40]
  wire [3:0] _GEN_467 = ~_GEN_127 ? _GEN_346 : _GEN_17; // @[ReservationStation.scala 66:40]
  wire [3:0] _GEN_468 = ~_GEN_127 ? _GEN_347 : _GEN_77; // @[ReservationStation.scala 66:40]
  wire [3:0] _GEN_469 = ~_GEN_127 ? _GEN_348 : _GEN_32; // @[ReservationStation.scala 66:40]
  wire [3:0] _GEN_470 = ~_GEN_127 ? _GEN_349 : _GEN_92; // @[ReservationStation.scala 66:40]
  wire [3:0] _GEN_471 = ~_GEN_127 ? _GEN_350 : _GEN_47; // @[ReservationStation.scala 66:40]
  wire [3:0] _GEN_472 = ~_GEN_127 ? _GEN_351 : _GEN_107; // @[ReservationStation.scala 66:40]
  wire  _GEN_473 = ~_GEN_127 ? _GEN_352 : _GEN_1; // @[ReservationStation.scala 66:40]
  wire  _GEN_474 = ~_GEN_127 ? _GEN_353 : _GEN_61; // @[ReservationStation.scala 66:40]
  wire  _GEN_475 = ~_GEN_127 ? _GEN_354 : _GEN_16; // @[ReservationStation.scala 66:40]
  wire  _GEN_476 = ~_GEN_127 ? _GEN_355 : _GEN_76; // @[ReservationStation.scala 66:40]
  wire  _GEN_477 = ~_GEN_127 ? _GEN_356 : _GEN_31; // @[ReservationStation.scala 66:40]
  wire  _GEN_478 = ~_GEN_127 ? _GEN_357 : _GEN_91; // @[ReservationStation.scala 66:40]
  wire  _GEN_479 = ~_GEN_127 ? _GEN_358 : _GEN_46; // @[ReservationStation.scala 66:40]
  wire  _GEN_480 = ~_GEN_127 ? _GEN_359 : _GEN_106; // @[ReservationStation.scala 66:40]
  wire  _GEN_481 = ~_GEN_127 ? _GEN_360 : _GEN_0; // @[ReservationStation.scala 66:40]
  wire  _GEN_482 = ~_GEN_127 ? _GEN_361 : _GEN_60; // @[ReservationStation.scala 66:40]
  wire  _GEN_483 = ~_GEN_127 ? _GEN_362 : _GEN_15; // @[ReservationStation.scala 66:40]
  wire  _GEN_484 = ~_GEN_127 ? _GEN_363 : _GEN_75; // @[ReservationStation.scala 66:40]
  wire  _GEN_485 = ~_GEN_127 ? _GEN_364 : _GEN_30; // @[ReservationStation.scala 66:40]
  wire  _GEN_486 = ~_GEN_127 ? _GEN_365 : _GEN_90; // @[ReservationStation.scala 66:40]
  wire  _GEN_487 = ~_GEN_127 ? _GEN_366 : _GEN_45; // @[ReservationStation.scala 66:40]
  wire  _GEN_488 = ~_GEN_127 ? _GEN_367 : _GEN_105; // @[ReservationStation.scala 66:40]
  wire  _T_10 = _T_8 & io_decoder_0_entry_valid; // @[ReservationStation.scala 73:36]
  wire [2:0] _T_12 = head + 3'h1; // @[ReservationStation.scala 74:16]
  wire [2:0] _T_13 = _T_10 ? _T_12 : head; // @[ReservationStation.scala 72:19]
  wire  _GEN_490 = 3'h1 == _T_13 ? reservation_1_valid : reservation_0_valid; // @[ReservationStation.scala 66:{10,10}]
  wire  _GEN_491 = 3'h2 == _T_13 ? reservation_2_valid : _GEN_490; // @[ReservationStation.scala 66:{10,10}]
  wire  _GEN_492 = 3'h3 == _T_13 ? reservation_3_valid : _GEN_491; // @[ReservationStation.scala 66:{10,10}]
  wire  _GEN_493 = 3'h4 == _T_13 ? reservation_4_valid : _GEN_492; // @[ReservationStation.scala 66:{10,10}]
  wire  _GEN_494 = 3'h5 == _T_13 ? reservation_5_valid : _GEN_493; // @[ReservationStation.scala 66:{10,10}]
  wire  _GEN_495 = 3'h6 == _T_13 ? reservation_6_valid : _GEN_494; // @[ReservationStation.scala 66:{10,10}]
  wire  _GEN_496 = 3'h7 == _T_13 ? reservation_7_valid : _GEN_495; // @[ReservationStation.scala 66:{10,10}]
  wire  _T_14 = ~_GEN_496; // @[ReservationStation.scala 66:10]
  wire  _GEN_537 = 3'h0 == _T_13 ? io_decoder_1_entry_ready1 : _GEN_409; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_538 = 3'h1 == _T_13 ? io_decoder_1_entry_ready1 : _GEN_410; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_539 = 3'h2 == _T_13 ? io_decoder_1_entry_ready1 : _GEN_411; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_540 = 3'h3 == _T_13 ? io_decoder_1_entry_ready1 : _GEN_412; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_541 = 3'h4 == _T_13 ? io_decoder_1_entry_ready1 : _GEN_413; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_542 = 3'h5 == _T_13 ? io_decoder_1_entry_ready1 : _GEN_414; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_543 = 3'h6 == _T_13 ? io_decoder_1_entry_ready1 : _GEN_415; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_544 = 3'h7 == _T_13 ? io_decoder_1_entry_ready1 : _GEN_416; // @[ReservationStation.scala 69:{31,31}]
  wire [63:0] _GEN_545 = 3'h0 == _T_13 ? io_decoder_1_entry_value1 : _GEN_417; // @[ReservationStation.scala 69:{31,31}]
  wire [63:0] _GEN_546 = 3'h1 == _T_13 ? io_decoder_1_entry_value1 : _GEN_418; // @[ReservationStation.scala 69:{31,31}]
  wire [63:0] _GEN_547 = 3'h2 == _T_13 ? io_decoder_1_entry_value1 : _GEN_419; // @[ReservationStation.scala 69:{31,31}]
  wire [63:0] _GEN_548 = 3'h3 == _T_13 ? io_decoder_1_entry_value1 : _GEN_420; // @[ReservationStation.scala 69:{31,31}]
  wire [63:0] _GEN_549 = 3'h4 == _T_13 ? io_decoder_1_entry_value1 : _GEN_421; // @[ReservationStation.scala 69:{31,31}]
  wire [63:0] _GEN_550 = 3'h5 == _T_13 ? io_decoder_1_entry_value1 : _GEN_422; // @[ReservationStation.scala 69:{31,31}]
  wire [63:0] _GEN_551 = 3'h6 == _T_13 ? io_decoder_1_entry_value1 : _GEN_423; // @[ReservationStation.scala 69:{31,31}]
  wire [63:0] _GEN_552 = 3'h7 == _T_13 ? io_decoder_1_entry_value1 : _GEN_424; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_569 = 3'h0 == _T_13 ? io_decoder_1_entry_ready2 : _GEN_441; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_570 = 3'h1 == _T_13 ? io_decoder_1_entry_ready2 : _GEN_442; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_571 = 3'h2 == _T_13 ? io_decoder_1_entry_ready2 : _GEN_443; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_572 = 3'h3 == _T_13 ? io_decoder_1_entry_ready2 : _GEN_444; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_573 = 3'h4 == _T_13 ? io_decoder_1_entry_ready2 : _GEN_445; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_574 = 3'h5 == _T_13 ? io_decoder_1_entry_ready2 : _GEN_446; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_575 = 3'h6 == _T_13 ? io_decoder_1_entry_ready2 : _GEN_447; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_576 = 3'h7 == _T_13 ? io_decoder_1_entry_ready2 : _GEN_448; // @[ReservationStation.scala 69:{31,31}]
  wire [63:0] _GEN_577 = 3'h0 == _T_13 ? io_decoder_1_entry_value2 : _GEN_449; // @[ReservationStation.scala 69:{31,31}]
  wire [63:0] _GEN_578 = 3'h1 == _T_13 ? io_decoder_1_entry_value2 : _GEN_450; // @[ReservationStation.scala 69:{31,31}]
  wire [63:0] _GEN_579 = 3'h2 == _T_13 ? io_decoder_1_entry_value2 : _GEN_451; // @[ReservationStation.scala 69:{31,31}]
  wire [63:0] _GEN_580 = 3'h3 == _T_13 ? io_decoder_1_entry_value2 : _GEN_452; // @[ReservationStation.scala 69:{31,31}]
  wire [63:0] _GEN_581 = 3'h4 == _T_13 ? io_decoder_1_entry_value2 : _GEN_453; // @[ReservationStation.scala 69:{31,31}]
  wire [63:0] _GEN_582 = 3'h5 == _T_13 ? io_decoder_1_entry_value2 : _GEN_454; // @[ReservationStation.scala 69:{31,31}]
  wire [63:0] _GEN_583 = 3'h6 == _T_13 ? io_decoder_1_entry_value2 : _GEN_455; // @[ReservationStation.scala 69:{31,31}]
  wire [63:0] _GEN_584 = 3'h7 == _T_13 ? io_decoder_1_entry_value2 : _GEN_456; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_585 = 3'h0 == _T_13 | _GEN_457; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_586 = 3'h1 == _T_13 | _GEN_458; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_587 = 3'h2 == _T_13 | _GEN_459; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_588 = 3'h3 == _T_13 | _GEN_460; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_589 = 3'h4 == _T_13 | _GEN_461; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_590 = 3'h5 == _T_13 | _GEN_462; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_591 = 3'h6 == _T_13 | _GEN_463; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_592 = 3'h7 == _T_13 | _GEN_464; // @[ReservationStation.scala 69:{31,31}]
  wire  _GEN_657 = io_decoder_1_entry_valid ? _GEN_537 : _GEN_409; // @[ReservationStation.scala 68:39]
  wire  _GEN_658 = io_decoder_1_entry_valid ? _GEN_538 : _GEN_410; // @[ReservationStation.scala 68:39]
  wire  _GEN_659 = io_decoder_1_entry_valid ? _GEN_539 : _GEN_411; // @[ReservationStation.scala 68:39]
  wire  _GEN_660 = io_decoder_1_entry_valid ? _GEN_540 : _GEN_412; // @[ReservationStation.scala 68:39]
  wire  _GEN_661 = io_decoder_1_entry_valid ? _GEN_541 : _GEN_413; // @[ReservationStation.scala 68:39]
  wire  _GEN_662 = io_decoder_1_entry_valid ? _GEN_542 : _GEN_414; // @[ReservationStation.scala 68:39]
  wire  _GEN_663 = io_decoder_1_entry_valid ? _GEN_543 : _GEN_415; // @[ReservationStation.scala 68:39]
  wire  _GEN_664 = io_decoder_1_entry_valid ? _GEN_544 : _GEN_416; // @[ReservationStation.scala 68:39]
  wire [63:0] _GEN_665 = io_decoder_1_entry_valid ? _GEN_545 : _GEN_417; // @[ReservationStation.scala 68:39]
  wire [63:0] _GEN_666 = io_decoder_1_entry_valid ? _GEN_546 : _GEN_418; // @[ReservationStation.scala 68:39]
  wire [63:0] _GEN_667 = io_decoder_1_entry_valid ? _GEN_547 : _GEN_419; // @[ReservationStation.scala 68:39]
  wire [63:0] _GEN_668 = io_decoder_1_entry_valid ? _GEN_548 : _GEN_420; // @[ReservationStation.scala 68:39]
  wire [63:0] _GEN_669 = io_decoder_1_entry_valid ? _GEN_549 : _GEN_421; // @[ReservationStation.scala 68:39]
  wire [63:0] _GEN_670 = io_decoder_1_entry_valid ? _GEN_550 : _GEN_422; // @[ReservationStation.scala 68:39]
  wire [63:0] _GEN_671 = io_decoder_1_entry_valid ? _GEN_551 : _GEN_423; // @[ReservationStation.scala 68:39]
  wire [63:0] _GEN_672 = io_decoder_1_entry_valid ? _GEN_552 : _GEN_424; // @[ReservationStation.scala 68:39]
  wire  _GEN_689 = io_decoder_1_entry_valid ? _GEN_569 : _GEN_441; // @[ReservationStation.scala 68:39]
  wire  _GEN_690 = io_decoder_1_entry_valid ? _GEN_570 : _GEN_442; // @[ReservationStation.scala 68:39]
  wire  _GEN_691 = io_decoder_1_entry_valid ? _GEN_571 : _GEN_443; // @[ReservationStation.scala 68:39]
  wire  _GEN_692 = io_decoder_1_entry_valid ? _GEN_572 : _GEN_444; // @[ReservationStation.scala 68:39]
  wire  _GEN_693 = io_decoder_1_entry_valid ? _GEN_573 : _GEN_445; // @[ReservationStation.scala 68:39]
  wire  _GEN_694 = io_decoder_1_entry_valid ? _GEN_574 : _GEN_446; // @[ReservationStation.scala 68:39]
  wire  _GEN_695 = io_decoder_1_entry_valid ? _GEN_575 : _GEN_447; // @[ReservationStation.scala 68:39]
  wire  _GEN_696 = io_decoder_1_entry_valid ? _GEN_576 : _GEN_448; // @[ReservationStation.scala 68:39]
  wire [63:0] _GEN_697 = io_decoder_1_entry_valid ? _GEN_577 : _GEN_449; // @[ReservationStation.scala 68:39]
  wire [63:0] _GEN_698 = io_decoder_1_entry_valid ? _GEN_578 : _GEN_450; // @[ReservationStation.scala 68:39]
  wire [63:0] _GEN_699 = io_decoder_1_entry_valid ? _GEN_579 : _GEN_451; // @[ReservationStation.scala 68:39]
  wire [63:0] _GEN_700 = io_decoder_1_entry_valid ? _GEN_580 : _GEN_452; // @[ReservationStation.scala 68:39]
  wire [63:0] _GEN_701 = io_decoder_1_entry_valid ? _GEN_581 : _GEN_453; // @[ReservationStation.scala 68:39]
  wire [63:0] _GEN_702 = io_decoder_1_entry_valid ? _GEN_582 : _GEN_454; // @[ReservationStation.scala 68:39]
  wire [63:0] _GEN_703 = io_decoder_1_entry_valid ? _GEN_583 : _GEN_455; // @[ReservationStation.scala 68:39]
  wire [63:0] _GEN_704 = io_decoder_1_entry_valid ? _GEN_584 : _GEN_456; // @[ReservationStation.scala 68:39]
  wire  _GEN_778 = ~_GEN_496 ? _GEN_657 : _GEN_409; // @[ReservationStation.scala 66:40]
  wire  _GEN_779 = ~_GEN_496 ? _GEN_658 : _GEN_410; // @[ReservationStation.scala 66:40]
  wire  _GEN_780 = ~_GEN_496 ? _GEN_659 : _GEN_411; // @[ReservationStation.scala 66:40]
  wire  _GEN_781 = ~_GEN_496 ? _GEN_660 : _GEN_412; // @[ReservationStation.scala 66:40]
  wire  _GEN_782 = ~_GEN_496 ? _GEN_661 : _GEN_413; // @[ReservationStation.scala 66:40]
  wire  _GEN_783 = ~_GEN_496 ? _GEN_662 : _GEN_414; // @[ReservationStation.scala 66:40]
  wire  _GEN_784 = ~_GEN_496 ? _GEN_663 : _GEN_415; // @[ReservationStation.scala 66:40]
  wire  _GEN_785 = ~_GEN_496 ? _GEN_664 : _GEN_416; // @[ReservationStation.scala 66:40]
  wire [63:0] _GEN_786 = ~_GEN_496 ? _GEN_665 : _GEN_417; // @[ReservationStation.scala 66:40]
  wire [63:0] _GEN_787 = ~_GEN_496 ? _GEN_666 : _GEN_418; // @[ReservationStation.scala 66:40]
  wire [63:0] _GEN_788 = ~_GEN_496 ? _GEN_667 : _GEN_419; // @[ReservationStation.scala 66:40]
  wire [63:0] _GEN_789 = ~_GEN_496 ? _GEN_668 : _GEN_420; // @[ReservationStation.scala 66:40]
  wire [63:0] _GEN_790 = ~_GEN_496 ? _GEN_669 : _GEN_421; // @[ReservationStation.scala 66:40]
  wire [63:0] _GEN_791 = ~_GEN_496 ? _GEN_670 : _GEN_422; // @[ReservationStation.scala 66:40]
  wire [63:0] _GEN_792 = ~_GEN_496 ? _GEN_671 : _GEN_423; // @[ReservationStation.scala 66:40]
  wire [63:0] _GEN_793 = ~_GEN_496 ? _GEN_672 : _GEN_424; // @[ReservationStation.scala 66:40]
  wire  _GEN_810 = ~_GEN_496 ? _GEN_689 : _GEN_441; // @[ReservationStation.scala 66:40]
  wire  _GEN_811 = ~_GEN_496 ? _GEN_690 : _GEN_442; // @[ReservationStation.scala 66:40]
  wire  _GEN_812 = ~_GEN_496 ? _GEN_691 : _GEN_443; // @[ReservationStation.scala 66:40]
  wire  _GEN_813 = ~_GEN_496 ? _GEN_692 : _GEN_444; // @[ReservationStation.scala 66:40]
  wire  _GEN_814 = ~_GEN_496 ? _GEN_693 : _GEN_445; // @[ReservationStation.scala 66:40]
  wire  _GEN_815 = ~_GEN_496 ? _GEN_694 : _GEN_446; // @[ReservationStation.scala 66:40]
  wire  _GEN_816 = ~_GEN_496 ? _GEN_695 : _GEN_447; // @[ReservationStation.scala 66:40]
  wire  _GEN_817 = ~_GEN_496 ? _GEN_696 : _GEN_448; // @[ReservationStation.scala 66:40]
  wire [63:0] _GEN_818 = ~_GEN_496 ? _GEN_697 : _GEN_449; // @[ReservationStation.scala 66:40]
  wire [63:0] _GEN_819 = ~_GEN_496 ? _GEN_698 : _GEN_450; // @[ReservationStation.scala 66:40]
  wire [63:0] _GEN_820 = ~_GEN_496 ? _GEN_699 : _GEN_451; // @[ReservationStation.scala 66:40]
  wire [63:0] _GEN_821 = ~_GEN_496 ? _GEN_700 : _GEN_452; // @[ReservationStation.scala 66:40]
  wire [63:0] _GEN_822 = ~_GEN_496 ? _GEN_701 : _GEN_453; // @[ReservationStation.scala 66:40]
  wire [63:0] _GEN_823 = ~_GEN_496 ? _GEN_702 : _GEN_454; // @[ReservationStation.scala 66:40]
  wire [63:0] _GEN_824 = ~_GEN_496 ? _GEN_703 : _GEN_455; // @[ReservationStation.scala 66:40]
  wire [63:0] _GEN_825 = ~_GEN_496 ? _GEN_704 : _GEN_456; // @[ReservationStation.scala 66:40]
  wire  _T_16 = _T_14 & io_decoder_1_entry_valid; // @[ReservationStation.scala 73:36]
  wire [2:0] _T_18 = _T_13 + 3'h1; // @[ReservationStation.scala 74:16]
  wire  _T_21 = io_collectedOutput_0_outputs_valid & ~io_collectedOutput_0_outputs_bits_resultType; // @[ReservationStation.scala 82:28]
  wire  _T_25 = reservation_0_sourceTag1_id == io_collectedOutput_0_outputs_bits_tag_id &
    reservation_0_sourceTag1_threadId == io_collectedOutput_0_outputs_bits_tag_threadId; // @[Tag.scala 13:25]
  wire [63:0] _GEN_858 = ~reservation_0_ready1 & _T_25 ? io_collectedOutput_0_outputs_bits_value : _GEN_786; // @[ReservationStation.scala 86:79 87:26]
  wire  _GEN_859 = ~reservation_0_ready1 & _T_25 | _GEN_778; // @[ReservationStation.scala 86:79 88:26]
  wire  _T_30 = reservation_0_sourceTag2_id == io_collectedOutput_0_outputs_bits_tag_id &
    reservation_0_sourceTag2_threadId == io_collectedOutput_0_outputs_bits_tag_threadId; // @[Tag.scala 13:25]
  wire [63:0] _GEN_860 = ~reservation_0_ready2 & _T_30 ? io_collectedOutput_0_outputs_bits_value : _GEN_818; // @[ReservationStation.scala 90:79 91:26]
  wire  _GEN_861 = ~reservation_0_ready2 & _T_30 | _GEN_810; // @[ReservationStation.scala 90:79 92:26]
  wire [63:0] _GEN_862 = reservation_0_valid ? _GEN_858 : _GEN_786; // @[ReservationStation.scala 85:27]
  wire  _GEN_863 = reservation_0_valid ? _GEN_859 : _GEN_778; // @[ReservationStation.scala 85:27]
  wire [63:0] _GEN_864 = reservation_0_valid ? _GEN_860 : _GEN_818; // @[ReservationStation.scala 85:27]
  wire  _GEN_865 = reservation_0_valid ? _GEN_861 : _GEN_810; // @[ReservationStation.scala 85:27]
  wire  _T_35 = reservation_1_sourceTag1_id == io_collectedOutput_0_outputs_bits_tag_id &
    reservation_1_sourceTag1_threadId == io_collectedOutput_0_outputs_bits_tag_threadId; // @[Tag.scala 13:25]
  wire [63:0] _GEN_866 = ~reservation_1_ready1 & _T_35 ? io_collectedOutput_0_outputs_bits_value : _GEN_787; // @[ReservationStation.scala 86:79 87:26]
  wire  _GEN_867 = ~reservation_1_ready1 & _T_35 | _GEN_779; // @[ReservationStation.scala 86:79 88:26]
  wire  _T_40 = reservation_1_sourceTag2_id == io_collectedOutput_0_outputs_bits_tag_id &
    reservation_1_sourceTag2_threadId == io_collectedOutput_0_outputs_bits_tag_threadId; // @[Tag.scala 13:25]
  wire [63:0] _GEN_868 = ~reservation_1_ready2 & _T_40 ? io_collectedOutput_0_outputs_bits_value : _GEN_819; // @[ReservationStation.scala 90:79 91:26]
  wire  _GEN_869 = ~reservation_1_ready2 & _T_40 | _GEN_811; // @[ReservationStation.scala 90:79 92:26]
  wire [63:0] _GEN_870 = reservation_1_valid ? _GEN_866 : _GEN_787; // @[ReservationStation.scala 85:27]
  wire  _GEN_871 = reservation_1_valid ? _GEN_867 : _GEN_779; // @[ReservationStation.scala 85:27]
  wire [63:0] _GEN_872 = reservation_1_valid ? _GEN_868 : _GEN_819; // @[ReservationStation.scala 85:27]
  wire  _GEN_873 = reservation_1_valid ? _GEN_869 : _GEN_811; // @[ReservationStation.scala 85:27]
  wire  _T_45 = reservation_2_sourceTag1_id == io_collectedOutput_0_outputs_bits_tag_id &
    reservation_2_sourceTag1_threadId == io_collectedOutput_0_outputs_bits_tag_threadId; // @[Tag.scala 13:25]
  wire [63:0] _GEN_874 = ~reservation_2_ready1 & _T_45 ? io_collectedOutput_0_outputs_bits_value : _GEN_788; // @[ReservationStation.scala 86:79 87:26]
  wire  _GEN_875 = ~reservation_2_ready1 & _T_45 | _GEN_780; // @[ReservationStation.scala 86:79 88:26]
  wire  _T_50 = reservation_2_sourceTag2_id == io_collectedOutput_0_outputs_bits_tag_id &
    reservation_2_sourceTag2_threadId == io_collectedOutput_0_outputs_bits_tag_threadId; // @[Tag.scala 13:25]
  wire [63:0] _GEN_876 = ~reservation_2_ready2 & _T_50 ? io_collectedOutput_0_outputs_bits_value : _GEN_820; // @[ReservationStation.scala 90:79 91:26]
  wire  _GEN_877 = ~reservation_2_ready2 & _T_50 | _GEN_812; // @[ReservationStation.scala 90:79 92:26]
  wire [63:0] _GEN_878 = reservation_2_valid ? _GEN_874 : _GEN_788; // @[ReservationStation.scala 85:27]
  wire  _GEN_879 = reservation_2_valid ? _GEN_875 : _GEN_780; // @[ReservationStation.scala 85:27]
  wire [63:0] _GEN_880 = reservation_2_valid ? _GEN_876 : _GEN_820; // @[ReservationStation.scala 85:27]
  wire  _GEN_881 = reservation_2_valid ? _GEN_877 : _GEN_812; // @[ReservationStation.scala 85:27]
  wire  _T_55 = reservation_3_sourceTag1_id == io_collectedOutput_0_outputs_bits_tag_id &
    reservation_3_sourceTag1_threadId == io_collectedOutput_0_outputs_bits_tag_threadId; // @[Tag.scala 13:25]
  wire [63:0] _GEN_882 = ~reservation_3_ready1 & _T_55 ? io_collectedOutput_0_outputs_bits_value : _GEN_789; // @[ReservationStation.scala 86:79 87:26]
  wire  _GEN_883 = ~reservation_3_ready1 & _T_55 | _GEN_781; // @[ReservationStation.scala 86:79 88:26]
  wire  _T_60 = reservation_3_sourceTag2_id == io_collectedOutput_0_outputs_bits_tag_id &
    reservation_3_sourceTag2_threadId == io_collectedOutput_0_outputs_bits_tag_threadId; // @[Tag.scala 13:25]
  wire [63:0] _GEN_884 = ~reservation_3_ready2 & _T_60 ? io_collectedOutput_0_outputs_bits_value : _GEN_821; // @[ReservationStation.scala 90:79 91:26]
  wire  _GEN_885 = ~reservation_3_ready2 & _T_60 | _GEN_813; // @[ReservationStation.scala 90:79 92:26]
  wire [63:0] _GEN_886 = reservation_3_valid ? _GEN_882 : _GEN_789; // @[ReservationStation.scala 85:27]
  wire  _GEN_887 = reservation_3_valid ? _GEN_883 : _GEN_781; // @[ReservationStation.scala 85:27]
  wire [63:0] _GEN_888 = reservation_3_valid ? _GEN_884 : _GEN_821; // @[ReservationStation.scala 85:27]
  wire  _GEN_889 = reservation_3_valid ? _GEN_885 : _GEN_813; // @[ReservationStation.scala 85:27]
  wire  _T_65 = reservation_4_sourceTag1_id == io_collectedOutput_0_outputs_bits_tag_id &
    reservation_4_sourceTag1_threadId == io_collectedOutput_0_outputs_bits_tag_threadId; // @[Tag.scala 13:25]
  wire [63:0] _GEN_890 = ~reservation_4_ready1 & _T_65 ? io_collectedOutput_0_outputs_bits_value : _GEN_790; // @[ReservationStation.scala 86:79 87:26]
  wire  _GEN_891 = ~reservation_4_ready1 & _T_65 | _GEN_782; // @[ReservationStation.scala 86:79 88:26]
  wire  _T_70 = reservation_4_sourceTag2_id == io_collectedOutput_0_outputs_bits_tag_id &
    reservation_4_sourceTag2_threadId == io_collectedOutput_0_outputs_bits_tag_threadId; // @[Tag.scala 13:25]
  wire [63:0] _GEN_892 = ~reservation_4_ready2 & _T_70 ? io_collectedOutput_0_outputs_bits_value : _GEN_822; // @[ReservationStation.scala 90:79 91:26]
  wire  _GEN_893 = ~reservation_4_ready2 & _T_70 | _GEN_814; // @[ReservationStation.scala 90:79 92:26]
  wire [63:0] _GEN_894 = reservation_4_valid ? _GEN_890 : _GEN_790; // @[ReservationStation.scala 85:27]
  wire  _GEN_895 = reservation_4_valid ? _GEN_891 : _GEN_782; // @[ReservationStation.scala 85:27]
  wire [63:0] _GEN_896 = reservation_4_valid ? _GEN_892 : _GEN_822; // @[ReservationStation.scala 85:27]
  wire  _GEN_897 = reservation_4_valid ? _GEN_893 : _GEN_814; // @[ReservationStation.scala 85:27]
  wire  _T_75 = reservation_5_sourceTag1_id == io_collectedOutput_0_outputs_bits_tag_id &
    reservation_5_sourceTag1_threadId == io_collectedOutput_0_outputs_bits_tag_threadId; // @[Tag.scala 13:25]
  wire [63:0] _GEN_898 = ~reservation_5_ready1 & _T_75 ? io_collectedOutput_0_outputs_bits_value : _GEN_791; // @[ReservationStation.scala 86:79 87:26]
  wire  _GEN_899 = ~reservation_5_ready1 & _T_75 | _GEN_783; // @[ReservationStation.scala 86:79 88:26]
  wire  _T_80 = reservation_5_sourceTag2_id == io_collectedOutput_0_outputs_bits_tag_id &
    reservation_5_sourceTag2_threadId == io_collectedOutput_0_outputs_bits_tag_threadId; // @[Tag.scala 13:25]
  wire [63:0] _GEN_900 = ~reservation_5_ready2 & _T_80 ? io_collectedOutput_0_outputs_bits_value : _GEN_823; // @[ReservationStation.scala 90:79 91:26]
  wire  _GEN_901 = ~reservation_5_ready2 & _T_80 | _GEN_815; // @[ReservationStation.scala 90:79 92:26]
  wire [63:0] _GEN_902 = reservation_5_valid ? _GEN_898 : _GEN_791; // @[ReservationStation.scala 85:27]
  wire  _GEN_903 = reservation_5_valid ? _GEN_899 : _GEN_783; // @[ReservationStation.scala 85:27]
  wire [63:0] _GEN_904 = reservation_5_valid ? _GEN_900 : _GEN_823; // @[ReservationStation.scala 85:27]
  wire  _GEN_905 = reservation_5_valid ? _GEN_901 : _GEN_815; // @[ReservationStation.scala 85:27]
  wire  _T_85 = reservation_6_sourceTag1_id == io_collectedOutput_0_outputs_bits_tag_id &
    reservation_6_sourceTag1_threadId == io_collectedOutput_0_outputs_bits_tag_threadId; // @[Tag.scala 13:25]
  wire [63:0] _GEN_906 = ~reservation_6_ready1 & _T_85 ? io_collectedOutput_0_outputs_bits_value : _GEN_792; // @[ReservationStation.scala 86:79 87:26]
  wire  _GEN_907 = ~reservation_6_ready1 & _T_85 | _GEN_784; // @[ReservationStation.scala 86:79 88:26]
  wire  _T_90 = reservation_6_sourceTag2_id == io_collectedOutput_0_outputs_bits_tag_id &
    reservation_6_sourceTag2_threadId == io_collectedOutput_0_outputs_bits_tag_threadId; // @[Tag.scala 13:25]
  wire [63:0] _GEN_908 = ~reservation_6_ready2 & _T_90 ? io_collectedOutput_0_outputs_bits_value : _GEN_824; // @[ReservationStation.scala 90:79 91:26]
  wire  _GEN_909 = ~reservation_6_ready2 & _T_90 | _GEN_816; // @[ReservationStation.scala 90:79 92:26]
  wire [63:0] _GEN_910 = reservation_6_valid ? _GEN_906 : _GEN_792; // @[ReservationStation.scala 85:27]
  wire  _GEN_911 = reservation_6_valid ? _GEN_907 : _GEN_784; // @[ReservationStation.scala 85:27]
  wire [63:0] _GEN_912 = reservation_6_valid ? _GEN_908 : _GEN_824; // @[ReservationStation.scala 85:27]
  wire  _GEN_913 = reservation_6_valid ? _GEN_909 : _GEN_816; // @[ReservationStation.scala 85:27]
  wire  _T_95 = reservation_7_sourceTag1_id == io_collectedOutput_0_outputs_bits_tag_id &
    reservation_7_sourceTag1_threadId == io_collectedOutput_0_outputs_bits_tag_threadId; // @[Tag.scala 13:25]
  wire [63:0] _GEN_914 = ~reservation_7_ready1 & _T_95 ? io_collectedOutput_0_outputs_bits_value : _GEN_793; // @[ReservationStation.scala 86:79 87:26]
  wire  _GEN_915 = ~reservation_7_ready1 & _T_95 | _GEN_785; // @[ReservationStation.scala 86:79 88:26]
  wire  _T_100 = reservation_7_sourceTag2_id == io_collectedOutput_0_outputs_bits_tag_id &
    reservation_7_sourceTag2_threadId == io_collectedOutput_0_outputs_bits_tag_threadId; // @[Tag.scala 13:25]
  wire [63:0] _GEN_916 = ~reservation_7_ready2 & _T_100 ? io_collectedOutput_0_outputs_bits_value : _GEN_825; // @[ReservationStation.scala 90:79 91:26]
  wire  _GEN_917 = ~reservation_7_ready2 & _T_100 | _GEN_817; // @[ReservationStation.scala 90:79 92:26]
  wire [63:0] _GEN_918 = reservation_7_valid ? _GEN_914 : _GEN_793; // @[ReservationStation.scala 85:27]
  wire  _GEN_919 = reservation_7_valid ? _GEN_915 : _GEN_785; // @[ReservationStation.scala 85:27]
  wire [63:0] _GEN_920 = reservation_7_valid ? _GEN_916 : _GEN_825; // @[ReservationStation.scala 85:27]
  wire  _GEN_921 = reservation_7_valid ? _GEN_917 : _GEN_817; // @[ReservationStation.scala 85:27]
  wire [63:0] _GEN_922 = _T_21 ? _GEN_862 : _GEN_786; // @[ReservationStation.scala 83:7]
  wire  _GEN_923 = _T_21 ? _GEN_863 : _GEN_778; // @[ReservationStation.scala 83:7]
  wire [63:0] _GEN_924 = _T_21 ? _GEN_864 : _GEN_818; // @[ReservationStation.scala 83:7]
  wire  _GEN_925 = _T_21 ? _GEN_865 : _GEN_810; // @[ReservationStation.scala 83:7]
  wire [63:0] _GEN_926 = _T_21 ? _GEN_870 : _GEN_787; // @[ReservationStation.scala 83:7]
  wire  _GEN_927 = _T_21 ? _GEN_871 : _GEN_779; // @[ReservationStation.scala 83:7]
  wire [63:0] _GEN_928 = _T_21 ? _GEN_872 : _GEN_819; // @[ReservationStation.scala 83:7]
  wire  _GEN_929 = _T_21 ? _GEN_873 : _GEN_811; // @[ReservationStation.scala 83:7]
  wire [63:0] _GEN_930 = _T_21 ? _GEN_878 : _GEN_788; // @[ReservationStation.scala 83:7]
  wire  _GEN_931 = _T_21 ? _GEN_879 : _GEN_780; // @[ReservationStation.scala 83:7]
  wire [63:0] _GEN_932 = _T_21 ? _GEN_880 : _GEN_820; // @[ReservationStation.scala 83:7]
  wire  _GEN_933 = _T_21 ? _GEN_881 : _GEN_812; // @[ReservationStation.scala 83:7]
  wire [63:0] _GEN_934 = _T_21 ? _GEN_886 : _GEN_789; // @[ReservationStation.scala 83:7]
  wire  _GEN_935 = _T_21 ? _GEN_887 : _GEN_781; // @[ReservationStation.scala 83:7]
  wire [63:0] _GEN_936 = _T_21 ? _GEN_888 : _GEN_821; // @[ReservationStation.scala 83:7]
  wire  _GEN_937 = _T_21 ? _GEN_889 : _GEN_813; // @[ReservationStation.scala 83:7]
  wire [63:0] _GEN_938 = _T_21 ? _GEN_894 : _GEN_790; // @[ReservationStation.scala 83:7]
  wire  _GEN_939 = _T_21 ? _GEN_895 : _GEN_782; // @[ReservationStation.scala 83:7]
  wire [63:0] _GEN_940 = _T_21 ? _GEN_896 : _GEN_822; // @[ReservationStation.scala 83:7]
  wire  _GEN_941 = _T_21 ? _GEN_897 : _GEN_814; // @[ReservationStation.scala 83:7]
  wire [63:0] _GEN_942 = _T_21 ? _GEN_902 : _GEN_791; // @[ReservationStation.scala 83:7]
  wire  _GEN_943 = _T_21 ? _GEN_903 : _GEN_783; // @[ReservationStation.scala 83:7]
  wire [63:0] _GEN_944 = _T_21 ? _GEN_904 : _GEN_823; // @[ReservationStation.scala 83:7]
  wire  _GEN_945 = _T_21 ? _GEN_905 : _GEN_815; // @[ReservationStation.scala 83:7]
  wire [63:0] _GEN_946 = _T_21 ? _GEN_910 : _GEN_792; // @[ReservationStation.scala 83:7]
  wire  _GEN_947 = _T_21 ? _GEN_911 : _GEN_784; // @[ReservationStation.scala 83:7]
  wire [63:0] _GEN_948 = _T_21 ? _GEN_912 : _GEN_824; // @[ReservationStation.scala 83:7]
  wire  _GEN_949 = _T_21 ? _GEN_913 : _GEN_816; // @[ReservationStation.scala 83:7]
  wire [63:0] _GEN_950 = _T_21 ? _GEN_918 : _GEN_793; // @[ReservationStation.scala 83:7]
  wire  _GEN_951 = _T_21 ? _GEN_919 : _GEN_785; // @[ReservationStation.scala 83:7]
  wire [63:0] _GEN_952 = _T_21 ? _GEN_920 : _GEN_825; // @[ReservationStation.scala 83:7]
  wire  _GEN_953 = _T_21 ? _GEN_921 : _GEN_817; // @[ReservationStation.scala 83:7]
  wire  _T_103 = io_collectedOutput_1_outputs_valid & ~io_collectedOutput_1_outputs_bits_resultType; // @[ReservationStation.scala 82:28]
  wire  _T_107 = reservation_0_sourceTag1_id == io_collectedOutput_1_outputs_bits_tag_id &
    reservation_0_sourceTag1_threadId == io_collectedOutput_1_outputs_bits_tag_threadId; // @[Tag.scala 13:25]
  wire  _GEN_955 = ~reservation_0_ready1 & _T_107 | _GEN_923; // @[ReservationStation.scala 86:79 88:26]
  wire  _T_112 = reservation_0_sourceTag2_id == io_collectedOutput_1_outputs_bits_tag_id &
    reservation_0_sourceTag2_threadId == io_collectedOutput_1_outputs_bits_tag_threadId; // @[Tag.scala 13:25]
  wire  _GEN_957 = ~reservation_0_ready2 & _T_112 | _GEN_925; // @[ReservationStation.scala 90:79 92:26]
  wire  _T_117 = reservation_1_sourceTag1_id == io_collectedOutput_1_outputs_bits_tag_id &
    reservation_1_sourceTag1_threadId == io_collectedOutput_1_outputs_bits_tag_threadId; // @[Tag.scala 13:25]
  wire  _GEN_963 = ~reservation_1_ready1 & _T_117 | _GEN_927; // @[ReservationStation.scala 86:79 88:26]
  wire  _T_122 = reservation_1_sourceTag2_id == io_collectedOutput_1_outputs_bits_tag_id &
    reservation_1_sourceTag2_threadId == io_collectedOutput_1_outputs_bits_tag_threadId; // @[Tag.scala 13:25]
  wire  _GEN_965 = ~reservation_1_ready2 & _T_122 | _GEN_929; // @[ReservationStation.scala 90:79 92:26]
  wire  _T_127 = reservation_2_sourceTag1_id == io_collectedOutput_1_outputs_bits_tag_id &
    reservation_2_sourceTag1_threadId == io_collectedOutput_1_outputs_bits_tag_threadId; // @[Tag.scala 13:25]
  wire  _GEN_971 = ~reservation_2_ready1 & _T_127 | _GEN_931; // @[ReservationStation.scala 86:79 88:26]
  wire  _T_132 = reservation_2_sourceTag2_id == io_collectedOutput_1_outputs_bits_tag_id &
    reservation_2_sourceTag2_threadId == io_collectedOutput_1_outputs_bits_tag_threadId; // @[Tag.scala 13:25]
  wire  _GEN_973 = ~reservation_2_ready2 & _T_132 | _GEN_933; // @[ReservationStation.scala 90:79 92:26]
  wire  _T_137 = reservation_3_sourceTag1_id == io_collectedOutput_1_outputs_bits_tag_id &
    reservation_3_sourceTag1_threadId == io_collectedOutput_1_outputs_bits_tag_threadId; // @[Tag.scala 13:25]
  wire  _GEN_979 = ~reservation_3_ready1 & _T_137 | _GEN_935; // @[ReservationStation.scala 86:79 88:26]
  wire  _T_142 = reservation_3_sourceTag2_id == io_collectedOutput_1_outputs_bits_tag_id &
    reservation_3_sourceTag2_threadId == io_collectedOutput_1_outputs_bits_tag_threadId; // @[Tag.scala 13:25]
  wire  _GEN_981 = ~reservation_3_ready2 & _T_142 | _GEN_937; // @[ReservationStation.scala 90:79 92:26]
  wire  _T_147 = reservation_4_sourceTag1_id == io_collectedOutput_1_outputs_bits_tag_id &
    reservation_4_sourceTag1_threadId == io_collectedOutput_1_outputs_bits_tag_threadId; // @[Tag.scala 13:25]
  wire  _GEN_987 = ~reservation_4_ready1 & _T_147 | _GEN_939; // @[ReservationStation.scala 86:79 88:26]
  wire  _T_152 = reservation_4_sourceTag2_id == io_collectedOutput_1_outputs_bits_tag_id &
    reservation_4_sourceTag2_threadId == io_collectedOutput_1_outputs_bits_tag_threadId; // @[Tag.scala 13:25]
  wire  _GEN_989 = ~reservation_4_ready2 & _T_152 | _GEN_941; // @[ReservationStation.scala 90:79 92:26]
  wire  _T_157 = reservation_5_sourceTag1_id == io_collectedOutput_1_outputs_bits_tag_id &
    reservation_5_sourceTag1_threadId == io_collectedOutput_1_outputs_bits_tag_threadId; // @[Tag.scala 13:25]
  wire  _GEN_995 = ~reservation_5_ready1 & _T_157 | _GEN_943; // @[ReservationStation.scala 86:79 88:26]
  wire  _T_162 = reservation_5_sourceTag2_id == io_collectedOutput_1_outputs_bits_tag_id &
    reservation_5_sourceTag2_threadId == io_collectedOutput_1_outputs_bits_tag_threadId; // @[Tag.scala 13:25]
  wire  _GEN_997 = ~reservation_5_ready2 & _T_162 | _GEN_945; // @[ReservationStation.scala 90:79 92:26]
  wire  _T_167 = reservation_6_sourceTag1_id == io_collectedOutput_1_outputs_bits_tag_id &
    reservation_6_sourceTag1_threadId == io_collectedOutput_1_outputs_bits_tag_threadId; // @[Tag.scala 13:25]
  wire  _GEN_1003 = ~reservation_6_ready1 & _T_167 | _GEN_947; // @[ReservationStation.scala 86:79 88:26]
  wire  _T_172 = reservation_6_sourceTag2_id == io_collectedOutput_1_outputs_bits_tag_id &
    reservation_6_sourceTag2_threadId == io_collectedOutput_1_outputs_bits_tag_threadId; // @[Tag.scala 13:25]
  wire  _GEN_1005 = ~reservation_6_ready2 & _T_172 | _GEN_949; // @[ReservationStation.scala 90:79 92:26]
  wire  _T_177 = reservation_7_sourceTag1_id == io_collectedOutput_1_outputs_bits_tag_id &
    reservation_7_sourceTag1_threadId == io_collectedOutput_1_outputs_bits_tag_threadId; // @[Tag.scala 13:25]
  wire  _GEN_1011 = ~reservation_7_ready1 & _T_177 | _GEN_951; // @[ReservationStation.scala 86:79 88:26]
  wire  _T_182 = reservation_7_sourceTag2_id == io_collectedOutput_1_outputs_bits_tag_id &
    reservation_7_sourceTag2_threadId == io_collectedOutput_1_outputs_bits_tag_threadId; // @[Tag.scala 13:25]
  wire  _GEN_1013 = ~reservation_7_ready2 & _T_182 | _GEN_953; // @[ReservationStation.scala 90:79 92:26]
  B4RRArbiter_1 outputArbiter_0 ( // @[ReservationStation.scala 34:11]
    .clock(outputArbiter_0_clock),
    .reset(outputArbiter_0_reset),
    .io_in_0_ready(outputArbiter_0_io_in_0_ready),
    .io_in_0_valid(outputArbiter_0_io_in_0_valid),
    .io_in_0_bits_destinationTag_threadId(outputArbiter_0_io_in_0_bits_destinationTag_threadId),
    .io_in_0_bits_destinationTag_id(outputArbiter_0_io_in_0_bits_destinationTag_id),
    .io_in_0_bits_value1(outputArbiter_0_io_in_0_bits_value1),
    .io_in_0_bits_value2(outputArbiter_0_io_in_0_bits_value2),
    .io_in_0_bits_function3(outputArbiter_0_io_in_0_bits_function3),
    .io_in_0_bits_immediateOrFunction7(outputArbiter_0_io_in_0_bits_immediateOrFunction7),
    .io_in_0_bits_opcode(outputArbiter_0_io_in_0_bits_opcode),
    .io_in_0_bits_wasCompressed(outputArbiter_0_io_in_0_bits_wasCompressed),
    .io_in_1_ready(outputArbiter_0_io_in_1_ready),
    .io_in_1_valid(outputArbiter_0_io_in_1_valid),
    .io_in_1_bits_destinationTag_threadId(outputArbiter_0_io_in_1_bits_destinationTag_threadId),
    .io_in_1_bits_destinationTag_id(outputArbiter_0_io_in_1_bits_destinationTag_id),
    .io_in_1_bits_value1(outputArbiter_0_io_in_1_bits_value1),
    .io_in_1_bits_value2(outputArbiter_0_io_in_1_bits_value2),
    .io_in_1_bits_function3(outputArbiter_0_io_in_1_bits_function3),
    .io_in_1_bits_immediateOrFunction7(outputArbiter_0_io_in_1_bits_immediateOrFunction7),
    .io_in_1_bits_opcode(outputArbiter_0_io_in_1_bits_opcode),
    .io_in_1_bits_wasCompressed(outputArbiter_0_io_in_1_bits_wasCompressed),
    .io_in_2_ready(outputArbiter_0_io_in_2_ready),
    .io_in_2_valid(outputArbiter_0_io_in_2_valid),
    .io_in_2_bits_destinationTag_threadId(outputArbiter_0_io_in_2_bits_destinationTag_threadId),
    .io_in_2_bits_destinationTag_id(outputArbiter_0_io_in_2_bits_destinationTag_id),
    .io_in_2_bits_value1(outputArbiter_0_io_in_2_bits_value1),
    .io_in_2_bits_value2(outputArbiter_0_io_in_2_bits_value2),
    .io_in_2_bits_function3(outputArbiter_0_io_in_2_bits_function3),
    .io_in_2_bits_immediateOrFunction7(outputArbiter_0_io_in_2_bits_immediateOrFunction7),
    .io_in_2_bits_opcode(outputArbiter_0_io_in_2_bits_opcode),
    .io_in_2_bits_wasCompressed(outputArbiter_0_io_in_2_bits_wasCompressed),
    .io_in_3_ready(outputArbiter_0_io_in_3_ready),
    .io_in_3_valid(outputArbiter_0_io_in_3_valid),
    .io_in_3_bits_destinationTag_threadId(outputArbiter_0_io_in_3_bits_destinationTag_threadId),
    .io_in_3_bits_destinationTag_id(outputArbiter_0_io_in_3_bits_destinationTag_id),
    .io_in_3_bits_value1(outputArbiter_0_io_in_3_bits_value1),
    .io_in_3_bits_value2(outputArbiter_0_io_in_3_bits_value2),
    .io_in_3_bits_function3(outputArbiter_0_io_in_3_bits_function3),
    .io_in_3_bits_immediateOrFunction7(outputArbiter_0_io_in_3_bits_immediateOrFunction7),
    .io_in_3_bits_opcode(outputArbiter_0_io_in_3_bits_opcode),
    .io_in_3_bits_wasCompressed(outputArbiter_0_io_in_3_bits_wasCompressed),
    .io_out_ready(outputArbiter_0_io_out_ready),
    .io_out_valid(outputArbiter_0_io_out_valid),
    .io_out_bits_destinationTag_threadId(outputArbiter_0_io_out_bits_destinationTag_threadId),
    .io_out_bits_destinationTag_id(outputArbiter_0_io_out_bits_destinationTag_id),
    .io_out_bits_value1(outputArbiter_0_io_out_bits_value1),
    .io_out_bits_value2(outputArbiter_0_io_out_bits_value2),
    .io_out_bits_function3(outputArbiter_0_io_out_bits_function3),
    .io_out_bits_immediateOrFunction7(outputArbiter_0_io_out_bits_immediateOrFunction7),
    .io_out_bits_opcode(outputArbiter_0_io_out_bits_opcode),
    .io_out_bits_wasCompressed(outputArbiter_0_io_out_bits_wasCompressed),
    .io_chosen(outputArbiter_0_io_chosen)
  );
  B4RRArbiter_1 outputArbiter_1 ( // @[ReservationStation.scala 34:11]
    .clock(outputArbiter_1_clock),
    .reset(outputArbiter_1_reset),
    .io_in_0_ready(outputArbiter_1_io_in_0_ready),
    .io_in_0_valid(outputArbiter_1_io_in_0_valid),
    .io_in_0_bits_destinationTag_threadId(outputArbiter_1_io_in_0_bits_destinationTag_threadId),
    .io_in_0_bits_destinationTag_id(outputArbiter_1_io_in_0_bits_destinationTag_id),
    .io_in_0_bits_value1(outputArbiter_1_io_in_0_bits_value1),
    .io_in_0_bits_value2(outputArbiter_1_io_in_0_bits_value2),
    .io_in_0_bits_function3(outputArbiter_1_io_in_0_bits_function3),
    .io_in_0_bits_immediateOrFunction7(outputArbiter_1_io_in_0_bits_immediateOrFunction7),
    .io_in_0_bits_opcode(outputArbiter_1_io_in_0_bits_opcode),
    .io_in_0_bits_wasCompressed(outputArbiter_1_io_in_0_bits_wasCompressed),
    .io_in_1_ready(outputArbiter_1_io_in_1_ready),
    .io_in_1_valid(outputArbiter_1_io_in_1_valid),
    .io_in_1_bits_destinationTag_threadId(outputArbiter_1_io_in_1_bits_destinationTag_threadId),
    .io_in_1_bits_destinationTag_id(outputArbiter_1_io_in_1_bits_destinationTag_id),
    .io_in_1_bits_value1(outputArbiter_1_io_in_1_bits_value1),
    .io_in_1_bits_value2(outputArbiter_1_io_in_1_bits_value2),
    .io_in_1_bits_function3(outputArbiter_1_io_in_1_bits_function3),
    .io_in_1_bits_immediateOrFunction7(outputArbiter_1_io_in_1_bits_immediateOrFunction7),
    .io_in_1_bits_opcode(outputArbiter_1_io_in_1_bits_opcode),
    .io_in_1_bits_wasCompressed(outputArbiter_1_io_in_1_bits_wasCompressed),
    .io_in_2_ready(outputArbiter_1_io_in_2_ready),
    .io_in_2_valid(outputArbiter_1_io_in_2_valid),
    .io_in_2_bits_destinationTag_threadId(outputArbiter_1_io_in_2_bits_destinationTag_threadId),
    .io_in_2_bits_destinationTag_id(outputArbiter_1_io_in_2_bits_destinationTag_id),
    .io_in_2_bits_value1(outputArbiter_1_io_in_2_bits_value1),
    .io_in_2_bits_value2(outputArbiter_1_io_in_2_bits_value2),
    .io_in_2_bits_function3(outputArbiter_1_io_in_2_bits_function3),
    .io_in_2_bits_immediateOrFunction7(outputArbiter_1_io_in_2_bits_immediateOrFunction7),
    .io_in_2_bits_opcode(outputArbiter_1_io_in_2_bits_opcode),
    .io_in_2_bits_wasCompressed(outputArbiter_1_io_in_2_bits_wasCompressed),
    .io_in_3_ready(outputArbiter_1_io_in_3_ready),
    .io_in_3_valid(outputArbiter_1_io_in_3_valid),
    .io_in_3_bits_destinationTag_threadId(outputArbiter_1_io_in_3_bits_destinationTag_threadId),
    .io_in_3_bits_destinationTag_id(outputArbiter_1_io_in_3_bits_destinationTag_id),
    .io_in_3_bits_value1(outputArbiter_1_io_in_3_bits_value1),
    .io_in_3_bits_value2(outputArbiter_1_io_in_3_bits_value2),
    .io_in_3_bits_function3(outputArbiter_1_io_in_3_bits_function3),
    .io_in_3_bits_immediateOrFunction7(outputArbiter_1_io_in_3_bits_immediateOrFunction7),
    .io_in_3_bits_opcode(outputArbiter_1_io_in_3_bits_opcode),
    .io_in_3_bits_wasCompressed(outputArbiter_1_io_in_3_bits_wasCompressed),
    .io_out_ready(outputArbiter_1_io_out_ready),
    .io_out_valid(outputArbiter_1_io_out_valid),
    .io_out_bits_destinationTag_threadId(outputArbiter_1_io_out_bits_destinationTag_threadId),
    .io_out_bits_destinationTag_id(outputArbiter_1_io_out_bits_destinationTag_id),
    .io_out_bits_value1(outputArbiter_1_io_out_bits_value1),
    .io_out_bits_value2(outputArbiter_1_io_out_bits_value2),
    .io_out_bits_function3(outputArbiter_1_io_out_bits_function3),
    .io_out_bits_immediateOrFunction7(outputArbiter_1_io_out_bits_immediateOrFunction7),
    .io_out_bits_opcode(outputArbiter_1_io_out_bits_opcode),
    .io_out_bits_wasCompressed(outputArbiter_1_io_out_bits_wasCompressed),
    .io_chosen(outputArbiter_1_io_chosen)
  );
  assign io_executor_0_valid = outputArbiter_0_io_out_valid; // @[ReservationStation.scala 58:22]
  assign io_executor_0_bits_destinationTag_threadId = outputArbiter_0_io_out_bits_destinationTag_threadId; // @[ReservationStation.scala 58:22]
  assign io_executor_0_bits_destinationTag_id = outputArbiter_0_io_out_bits_destinationTag_id; // @[ReservationStation.scala 58:22]
  assign io_executor_0_bits_value1 = outputArbiter_0_io_out_bits_value1; // @[ReservationStation.scala 58:22]
  assign io_executor_0_bits_value2 = outputArbiter_0_io_out_bits_value2; // @[ReservationStation.scala 58:22]
  assign io_executor_0_bits_function3 = outputArbiter_0_io_out_bits_function3; // @[ReservationStation.scala 58:22]
  assign io_executor_0_bits_immediateOrFunction7 = outputArbiter_0_io_out_bits_immediateOrFunction7; // @[ReservationStation.scala 58:22]
  assign io_executor_0_bits_opcode = outputArbiter_0_io_out_bits_opcode; // @[ReservationStation.scala 58:22]
  assign io_executor_0_bits_wasCompressed = outputArbiter_0_io_out_bits_wasCompressed; // @[ReservationStation.scala 58:22]
  assign io_executor_1_valid = outputArbiter_1_io_out_valid; // @[ReservationStation.scala 58:22]
  assign io_executor_1_bits_destinationTag_threadId = outputArbiter_1_io_out_bits_destinationTag_threadId; // @[ReservationStation.scala 58:22]
  assign io_executor_1_bits_destinationTag_id = outputArbiter_1_io_out_bits_destinationTag_id; // @[ReservationStation.scala 58:22]
  assign io_executor_1_bits_value1 = outputArbiter_1_io_out_bits_value1; // @[ReservationStation.scala 58:22]
  assign io_executor_1_bits_value2 = outputArbiter_1_io_out_bits_value2; // @[ReservationStation.scala 58:22]
  assign io_executor_1_bits_function3 = outputArbiter_1_io_out_bits_function3; // @[ReservationStation.scala 58:22]
  assign io_executor_1_bits_immediateOrFunction7 = outputArbiter_1_io_out_bits_immediateOrFunction7; // @[ReservationStation.scala 58:22]
  assign io_executor_1_bits_opcode = outputArbiter_1_io_out_bits_opcode; // @[ReservationStation.scala 58:22]
  assign io_executor_1_bits_wasCompressed = outputArbiter_1_io_out_bits_wasCompressed; // @[ReservationStation.scala 58:22]
  assign io_decoder_0_ready = ~_GEN_127; // @[ReservationStation.scala 66:10]
  assign io_decoder_1_ready = ~_GEN_496; // @[ReservationStation.scala 66:10]
  assign outputArbiter_0_clock = clock;
  assign outputArbiter_0_reset = reset;
  assign outputArbiter_0_io_in_0_valid = reservation_0_ready1 & reservation_0_ready2; // @[ReservationStation.scala 53:27]
  assign outputArbiter_0_io_in_0_bits_destinationTag_threadId = reservation_0_destinationTag_threadId; // @[ReservationStation.scala 47:29]
  assign outputArbiter_0_io_in_0_bits_destinationTag_id = reservation_0_destinationTag_id; // @[ReservationStation.scala 47:29]
  assign outputArbiter_0_io_in_0_bits_value1 = reservation_0_value1; // @[ReservationStation.scala 48:21]
  assign outputArbiter_0_io_in_0_bits_value2 = reservation_0_value2; // @[ReservationStation.scala 49:21]
  assign outputArbiter_0_io_in_0_bits_function3 = reservation_0_function3; // @[ReservationStation.scala 50:24]
  assign outputArbiter_0_io_in_0_bits_immediateOrFunction7 = reservation_0_immediateOrFunction7; // @[ReservationStation.scala 51:35]
  assign outputArbiter_0_io_in_0_bits_opcode = reservation_0_opcode; // @[ReservationStation.scala 46:21]
  assign outputArbiter_0_io_in_0_bits_wasCompressed = reservation_0_wasCompressed; // @[ReservationStation.scala 52:28]
  assign outputArbiter_0_io_in_1_valid = reservation_2_ready1 & reservation_2_ready2; // @[ReservationStation.scala 53:27]
  assign outputArbiter_0_io_in_1_bits_destinationTag_threadId = reservation_2_destinationTag_threadId; // @[ReservationStation.scala 47:29]
  assign outputArbiter_0_io_in_1_bits_destinationTag_id = reservation_2_destinationTag_id; // @[ReservationStation.scala 47:29]
  assign outputArbiter_0_io_in_1_bits_value1 = reservation_2_value1; // @[ReservationStation.scala 48:21]
  assign outputArbiter_0_io_in_1_bits_value2 = reservation_2_value2; // @[ReservationStation.scala 49:21]
  assign outputArbiter_0_io_in_1_bits_function3 = reservation_2_function3; // @[ReservationStation.scala 50:24]
  assign outputArbiter_0_io_in_1_bits_immediateOrFunction7 = reservation_2_immediateOrFunction7; // @[ReservationStation.scala 51:35]
  assign outputArbiter_0_io_in_1_bits_opcode = reservation_2_opcode; // @[ReservationStation.scala 46:21]
  assign outputArbiter_0_io_in_1_bits_wasCompressed = reservation_2_wasCompressed; // @[ReservationStation.scala 52:28]
  assign outputArbiter_0_io_in_2_valid = reservation_4_ready1 & reservation_4_ready2; // @[ReservationStation.scala 53:27]
  assign outputArbiter_0_io_in_2_bits_destinationTag_threadId = reservation_4_destinationTag_threadId; // @[ReservationStation.scala 47:29]
  assign outputArbiter_0_io_in_2_bits_destinationTag_id = reservation_4_destinationTag_id; // @[ReservationStation.scala 47:29]
  assign outputArbiter_0_io_in_2_bits_value1 = reservation_4_value1; // @[ReservationStation.scala 48:21]
  assign outputArbiter_0_io_in_2_bits_value2 = reservation_4_value2; // @[ReservationStation.scala 49:21]
  assign outputArbiter_0_io_in_2_bits_function3 = reservation_4_function3; // @[ReservationStation.scala 50:24]
  assign outputArbiter_0_io_in_2_bits_immediateOrFunction7 = reservation_4_immediateOrFunction7; // @[ReservationStation.scala 51:35]
  assign outputArbiter_0_io_in_2_bits_opcode = reservation_4_opcode; // @[ReservationStation.scala 46:21]
  assign outputArbiter_0_io_in_2_bits_wasCompressed = reservation_4_wasCompressed; // @[ReservationStation.scala 52:28]
  assign outputArbiter_0_io_in_3_valid = reservation_6_ready1 & reservation_6_ready2; // @[ReservationStation.scala 53:27]
  assign outputArbiter_0_io_in_3_bits_destinationTag_threadId = reservation_6_destinationTag_threadId; // @[ReservationStation.scala 47:29]
  assign outputArbiter_0_io_in_3_bits_destinationTag_id = reservation_6_destinationTag_id; // @[ReservationStation.scala 47:29]
  assign outputArbiter_0_io_in_3_bits_value1 = reservation_6_value1; // @[ReservationStation.scala 48:21]
  assign outputArbiter_0_io_in_3_bits_value2 = reservation_6_value2; // @[ReservationStation.scala 49:21]
  assign outputArbiter_0_io_in_3_bits_function3 = reservation_6_function3; // @[ReservationStation.scala 50:24]
  assign outputArbiter_0_io_in_3_bits_immediateOrFunction7 = reservation_6_immediateOrFunction7; // @[ReservationStation.scala 51:35]
  assign outputArbiter_0_io_in_3_bits_opcode = reservation_6_opcode; // @[ReservationStation.scala 46:21]
  assign outputArbiter_0_io_in_3_bits_wasCompressed = reservation_6_wasCompressed; // @[ReservationStation.scala 52:28]
  assign outputArbiter_0_io_out_ready = io_executor_0_ready; // @[ReservationStation.scala 58:22]
  assign outputArbiter_1_clock = clock;
  assign outputArbiter_1_reset = reset;
  assign outputArbiter_1_io_in_0_valid = reservation_1_ready1 & reservation_1_ready2; // @[ReservationStation.scala 53:27]
  assign outputArbiter_1_io_in_0_bits_destinationTag_threadId = reservation_1_destinationTag_threadId; // @[ReservationStation.scala 47:29]
  assign outputArbiter_1_io_in_0_bits_destinationTag_id = reservation_1_destinationTag_id; // @[ReservationStation.scala 47:29]
  assign outputArbiter_1_io_in_0_bits_value1 = reservation_1_value1; // @[ReservationStation.scala 48:21]
  assign outputArbiter_1_io_in_0_bits_value2 = reservation_1_value2; // @[ReservationStation.scala 49:21]
  assign outputArbiter_1_io_in_0_bits_function3 = reservation_1_function3; // @[ReservationStation.scala 50:24]
  assign outputArbiter_1_io_in_0_bits_immediateOrFunction7 = reservation_1_immediateOrFunction7; // @[ReservationStation.scala 51:35]
  assign outputArbiter_1_io_in_0_bits_opcode = reservation_1_opcode; // @[ReservationStation.scala 46:21]
  assign outputArbiter_1_io_in_0_bits_wasCompressed = reservation_1_wasCompressed; // @[ReservationStation.scala 52:28]
  assign outputArbiter_1_io_in_1_valid = reservation_3_ready1 & reservation_3_ready2; // @[ReservationStation.scala 53:27]
  assign outputArbiter_1_io_in_1_bits_destinationTag_threadId = reservation_3_destinationTag_threadId; // @[ReservationStation.scala 47:29]
  assign outputArbiter_1_io_in_1_bits_destinationTag_id = reservation_3_destinationTag_id; // @[ReservationStation.scala 47:29]
  assign outputArbiter_1_io_in_1_bits_value1 = reservation_3_value1; // @[ReservationStation.scala 48:21]
  assign outputArbiter_1_io_in_1_bits_value2 = reservation_3_value2; // @[ReservationStation.scala 49:21]
  assign outputArbiter_1_io_in_1_bits_function3 = reservation_3_function3; // @[ReservationStation.scala 50:24]
  assign outputArbiter_1_io_in_1_bits_immediateOrFunction7 = reservation_3_immediateOrFunction7; // @[ReservationStation.scala 51:35]
  assign outputArbiter_1_io_in_1_bits_opcode = reservation_3_opcode; // @[ReservationStation.scala 46:21]
  assign outputArbiter_1_io_in_1_bits_wasCompressed = reservation_3_wasCompressed; // @[ReservationStation.scala 52:28]
  assign outputArbiter_1_io_in_2_valid = reservation_5_ready1 & reservation_5_ready2; // @[ReservationStation.scala 53:27]
  assign outputArbiter_1_io_in_2_bits_destinationTag_threadId = reservation_5_destinationTag_threadId; // @[ReservationStation.scala 47:29]
  assign outputArbiter_1_io_in_2_bits_destinationTag_id = reservation_5_destinationTag_id; // @[ReservationStation.scala 47:29]
  assign outputArbiter_1_io_in_2_bits_value1 = reservation_5_value1; // @[ReservationStation.scala 48:21]
  assign outputArbiter_1_io_in_2_bits_value2 = reservation_5_value2; // @[ReservationStation.scala 49:21]
  assign outputArbiter_1_io_in_2_bits_function3 = reservation_5_function3; // @[ReservationStation.scala 50:24]
  assign outputArbiter_1_io_in_2_bits_immediateOrFunction7 = reservation_5_immediateOrFunction7; // @[ReservationStation.scala 51:35]
  assign outputArbiter_1_io_in_2_bits_opcode = reservation_5_opcode; // @[ReservationStation.scala 46:21]
  assign outputArbiter_1_io_in_2_bits_wasCompressed = reservation_5_wasCompressed; // @[ReservationStation.scala 52:28]
  assign outputArbiter_1_io_in_3_valid = reservation_7_ready1 & reservation_7_ready2; // @[ReservationStation.scala 53:27]
  assign outputArbiter_1_io_in_3_bits_destinationTag_threadId = reservation_7_destinationTag_threadId; // @[ReservationStation.scala 47:29]
  assign outputArbiter_1_io_in_3_bits_destinationTag_id = reservation_7_destinationTag_id; // @[ReservationStation.scala 47:29]
  assign outputArbiter_1_io_in_3_bits_value1 = reservation_7_value1; // @[ReservationStation.scala 48:21]
  assign outputArbiter_1_io_in_3_bits_value2 = reservation_7_value2; // @[ReservationStation.scala 49:21]
  assign outputArbiter_1_io_in_3_bits_function3 = reservation_7_function3; // @[ReservationStation.scala 50:24]
  assign outputArbiter_1_io_in_3_bits_immediateOrFunction7 = reservation_7_immediateOrFunction7; // @[ReservationStation.scala 51:35]
  assign outputArbiter_1_io_in_3_bits_opcode = reservation_7_opcode; // @[ReservationStation.scala 46:21]
  assign outputArbiter_1_io_in_3_bits_wasCompressed = reservation_7_wasCompressed; // @[ReservationStation.scala 52:28]
  assign outputArbiter_1_io_out_ready = io_executor_1_ready; // @[ReservationStation.scala 58:22]
  always @(posedge clock) begin
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_0_opcode <= 7'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h0 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_0_opcode <= io_decoder_1_entry_opcode; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_0_opcode <= _GEN_369;
        end
      end else begin
        reservation_0_opcode <= _GEN_369;
      end
    end else begin
      reservation_0_opcode <= _GEN_369;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_0_function3 <= 3'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h0 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_0_function3 <= io_decoder_1_entry_function3; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_0_function3 <= _GEN_377;
        end
      end else begin
        reservation_0_function3 <= _GEN_377;
      end
    end else begin
      reservation_0_function3 <= _GEN_377;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_0_immediateOrFunction7 <= 12'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h0 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_0_immediateOrFunction7 <= io_decoder_1_entry_immediateOrFunction7; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_0_immediateOrFunction7 <= _GEN_385;
        end
      end else begin
        reservation_0_immediateOrFunction7 <= _GEN_385;
      end
    end else begin
      reservation_0_immediateOrFunction7 <= _GEN_385;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_0_sourceTag1_threadId <= 1'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h0 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_0_sourceTag1_threadId <= io_decoder_1_entry_sourceTag1_threadId; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_0_sourceTag1_threadId <= _GEN_393;
        end
      end else begin
        reservation_0_sourceTag1_threadId <= _GEN_393;
      end
    end else begin
      reservation_0_sourceTag1_threadId <= _GEN_393;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_0_sourceTag1_id <= 4'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h0 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_0_sourceTag1_id <= io_decoder_1_entry_sourceTag1_id; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_0_sourceTag1_id <= _GEN_401;
        end
      end else begin
        reservation_0_sourceTag1_id <= _GEN_401;
      end
    end else begin
      reservation_0_sourceTag1_id <= _GEN_401;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_0_ready1 <= 1'h0; // @[ReservationStation.scala 28:28]
    end else if (_T_103) begin // @[ReservationStation.scala 83:7]
      if (reservation_0_valid) begin // @[ReservationStation.scala 85:27]
        reservation_0_ready1 <= _GEN_955;
      end else begin
        reservation_0_ready1 <= _GEN_923;
      end
    end else begin
      reservation_0_ready1 <= _GEN_923;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_0_value1 <= 64'h0; // @[ReservationStation.scala 28:28]
    end else if (_T_103) begin // @[ReservationStation.scala 83:7]
      if (reservation_0_valid) begin // @[ReservationStation.scala 85:27]
        if (~reservation_0_ready1 & _T_107) begin // @[ReservationStation.scala 86:79]
          reservation_0_value1 <= io_collectedOutput_1_outputs_bits_value; // @[ReservationStation.scala 87:26]
        end else begin
          reservation_0_value1 <= _GEN_922;
        end
      end else begin
        reservation_0_value1 <= _GEN_922;
      end
    end else begin
      reservation_0_value1 <= _GEN_922;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_0_sourceTag2_threadId <= 1'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h0 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_0_sourceTag2_threadId <= io_decoder_1_entry_sourceTag2_threadId; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_0_sourceTag2_threadId <= _GEN_425;
        end
      end else begin
        reservation_0_sourceTag2_threadId <= _GEN_425;
      end
    end else begin
      reservation_0_sourceTag2_threadId <= _GEN_425;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_0_sourceTag2_id <= 4'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h0 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_0_sourceTag2_id <= io_decoder_1_entry_sourceTag2_id; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_0_sourceTag2_id <= _GEN_433;
        end
      end else begin
        reservation_0_sourceTag2_id <= _GEN_433;
      end
    end else begin
      reservation_0_sourceTag2_id <= _GEN_433;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_0_ready2 <= 1'h0; // @[ReservationStation.scala 28:28]
    end else if (_T_103) begin // @[ReservationStation.scala 83:7]
      if (reservation_0_valid) begin // @[ReservationStation.scala 85:27]
        reservation_0_ready2 <= _GEN_957;
      end else begin
        reservation_0_ready2 <= _GEN_925;
      end
    end else begin
      reservation_0_ready2 <= _GEN_925;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_0_value2 <= 64'h0; // @[ReservationStation.scala 28:28]
    end else if (_T_103) begin // @[ReservationStation.scala 83:7]
      if (reservation_0_valid) begin // @[ReservationStation.scala 85:27]
        if (~reservation_0_ready2 & _T_112) begin // @[ReservationStation.scala 90:79]
          reservation_0_value2 <= io_collectedOutput_1_outputs_bits_value; // @[ReservationStation.scala 91:26]
        end else begin
          reservation_0_value2 <= _GEN_924;
        end
      end else begin
        reservation_0_value2 <= _GEN_924;
      end
    end else begin
      reservation_0_value2 <= _GEN_924;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_0_destinationTag_threadId <= 1'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        reservation_0_destinationTag_threadId <= _GEN_585;
      end else begin
        reservation_0_destinationTag_threadId <= _GEN_457;
      end
    end else begin
      reservation_0_destinationTag_threadId <= _GEN_457;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_0_destinationTag_id <= 4'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h0 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_0_destinationTag_id <= io_decoder_1_entry_destinationTag_id; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_0_destinationTag_id <= _GEN_465;
        end
      end else begin
        reservation_0_destinationTag_id <= _GEN_465;
      end
    end else begin
      reservation_0_destinationTag_id <= _GEN_465;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_0_wasCompressed <= 1'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h0 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_0_wasCompressed <= io_decoder_1_entry_wasCompressed; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_0_wasCompressed <= _GEN_473;
        end
      end else begin
        reservation_0_wasCompressed <= _GEN_473;
      end
    end else begin
      reservation_0_wasCompressed <= _GEN_473;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_0_valid <= 1'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h0 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_0_valid <= io_decoder_1_entry_valid; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_0_valid <= _GEN_481;
        end
      end else begin
        reservation_0_valid <= _GEN_481;
      end
    end else begin
      reservation_0_valid <= _GEN_481;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_1_opcode <= 7'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h1 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_1_opcode <= io_decoder_1_entry_opcode; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_1_opcode <= _GEN_370;
        end
      end else begin
        reservation_1_opcode <= _GEN_370;
      end
    end else begin
      reservation_1_opcode <= _GEN_370;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_1_function3 <= 3'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h1 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_1_function3 <= io_decoder_1_entry_function3; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_1_function3 <= _GEN_378;
        end
      end else begin
        reservation_1_function3 <= _GEN_378;
      end
    end else begin
      reservation_1_function3 <= _GEN_378;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_1_immediateOrFunction7 <= 12'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h1 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_1_immediateOrFunction7 <= io_decoder_1_entry_immediateOrFunction7; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_1_immediateOrFunction7 <= _GEN_386;
        end
      end else begin
        reservation_1_immediateOrFunction7 <= _GEN_386;
      end
    end else begin
      reservation_1_immediateOrFunction7 <= _GEN_386;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_1_sourceTag1_threadId <= 1'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h1 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_1_sourceTag1_threadId <= io_decoder_1_entry_sourceTag1_threadId; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_1_sourceTag1_threadId <= _GEN_394;
        end
      end else begin
        reservation_1_sourceTag1_threadId <= _GEN_394;
      end
    end else begin
      reservation_1_sourceTag1_threadId <= _GEN_394;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_1_sourceTag1_id <= 4'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h1 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_1_sourceTag1_id <= io_decoder_1_entry_sourceTag1_id; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_1_sourceTag1_id <= _GEN_402;
        end
      end else begin
        reservation_1_sourceTag1_id <= _GEN_402;
      end
    end else begin
      reservation_1_sourceTag1_id <= _GEN_402;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_1_ready1 <= 1'h0; // @[ReservationStation.scala 28:28]
    end else if (_T_103) begin // @[ReservationStation.scala 83:7]
      if (reservation_1_valid) begin // @[ReservationStation.scala 85:27]
        reservation_1_ready1 <= _GEN_963;
      end else begin
        reservation_1_ready1 <= _GEN_927;
      end
    end else begin
      reservation_1_ready1 <= _GEN_927;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_1_value1 <= 64'h0; // @[ReservationStation.scala 28:28]
    end else if (_T_103) begin // @[ReservationStation.scala 83:7]
      if (reservation_1_valid) begin // @[ReservationStation.scala 85:27]
        if (~reservation_1_ready1 & _T_117) begin // @[ReservationStation.scala 86:79]
          reservation_1_value1 <= io_collectedOutput_1_outputs_bits_value; // @[ReservationStation.scala 87:26]
        end else begin
          reservation_1_value1 <= _GEN_926;
        end
      end else begin
        reservation_1_value1 <= _GEN_926;
      end
    end else begin
      reservation_1_value1 <= _GEN_926;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_1_sourceTag2_threadId <= 1'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h1 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_1_sourceTag2_threadId <= io_decoder_1_entry_sourceTag2_threadId; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_1_sourceTag2_threadId <= _GEN_426;
        end
      end else begin
        reservation_1_sourceTag2_threadId <= _GEN_426;
      end
    end else begin
      reservation_1_sourceTag2_threadId <= _GEN_426;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_1_sourceTag2_id <= 4'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h1 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_1_sourceTag2_id <= io_decoder_1_entry_sourceTag2_id; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_1_sourceTag2_id <= _GEN_434;
        end
      end else begin
        reservation_1_sourceTag2_id <= _GEN_434;
      end
    end else begin
      reservation_1_sourceTag2_id <= _GEN_434;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_1_ready2 <= 1'h0; // @[ReservationStation.scala 28:28]
    end else if (_T_103) begin // @[ReservationStation.scala 83:7]
      if (reservation_1_valid) begin // @[ReservationStation.scala 85:27]
        reservation_1_ready2 <= _GEN_965;
      end else begin
        reservation_1_ready2 <= _GEN_929;
      end
    end else begin
      reservation_1_ready2 <= _GEN_929;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_1_value2 <= 64'h0; // @[ReservationStation.scala 28:28]
    end else if (_T_103) begin // @[ReservationStation.scala 83:7]
      if (reservation_1_valid) begin // @[ReservationStation.scala 85:27]
        if (~reservation_1_ready2 & _T_122) begin // @[ReservationStation.scala 90:79]
          reservation_1_value2 <= io_collectedOutput_1_outputs_bits_value; // @[ReservationStation.scala 91:26]
        end else begin
          reservation_1_value2 <= _GEN_928;
        end
      end else begin
        reservation_1_value2 <= _GEN_928;
      end
    end else begin
      reservation_1_value2 <= _GEN_928;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_1_destinationTag_threadId <= 1'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        reservation_1_destinationTag_threadId <= _GEN_586;
      end else begin
        reservation_1_destinationTag_threadId <= _GEN_458;
      end
    end else begin
      reservation_1_destinationTag_threadId <= _GEN_458;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_1_destinationTag_id <= 4'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h1 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_1_destinationTag_id <= io_decoder_1_entry_destinationTag_id; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_1_destinationTag_id <= _GEN_466;
        end
      end else begin
        reservation_1_destinationTag_id <= _GEN_466;
      end
    end else begin
      reservation_1_destinationTag_id <= _GEN_466;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_1_wasCompressed <= 1'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h1 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_1_wasCompressed <= io_decoder_1_entry_wasCompressed; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_1_wasCompressed <= _GEN_474;
        end
      end else begin
        reservation_1_wasCompressed <= _GEN_474;
      end
    end else begin
      reservation_1_wasCompressed <= _GEN_474;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_1_valid <= 1'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h1 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_1_valid <= io_decoder_1_entry_valid; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_1_valid <= _GEN_482;
        end
      end else begin
        reservation_1_valid <= _GEN_482;
      end
    end else begin
      reservation_1_valid <= _GEN_482;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_2_opcode <= 7'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h2 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_2_opcode <= io_decoder_1_entry_opcode; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_2_opcode <= _GEN_371;
        end
      end else begin
        reservation_2_opcode <= _GEN_371;
      end
    end else begin
      reservation_2_opcode <= _GEN_371;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_2_function3 <= 3'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h2 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_2_function3 <= io_decoder_1_entry_function3; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_2_function3 <= _GEN_379;
        end
      end else begin
        reservation_2_function3 <= _GEN_379;
      end
    end else begin
      reservation_2_function3 <= _GEN_379;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_2_immediateOrFunction7 <= 12'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h2 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_2_immediateOrFunction7 <= io_decoder_1_entry_immediateOrFunction7; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_2_immediateOrFunction7 <= _GEN_387;
        end
      end else begin
        reservation_2_immediateOrFunction7 <= _GEN_387;
      end
    end else begin
      reservation_2_immediateOrFunction7 <= _GEN_387;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_2_sourceTag1_threadId <= 1'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h2 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_2_sourceTag1_threadId <= io_decoder_1_entry_sourceTag1_threadId; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_2_sourceTag1_threadId <= _GEN_395;
        end
      end else begin
        reservation_2_sourceTag1_threadId <= _GEN_395;
      end
    end else begin
      reservation_2_sourceTag1_threadId <= _GEN_395;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_2_sourceTag1_id <= 4'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h2 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_2_sourceTag1_id <= io_decoder_1_entry_sourceTag1_id; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_2_sourceTag1_id <= _GEN_403;
        end
      end else begin
        reservation_2_sourceTag1_id <= _GEN_403;
      end
    end else begin
      reservation_2_sourceTag1_id <= _GEN_403;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_2_ready1 <= 1'h0; // @[ReservationStation.scala 28:28]
    end else if (_T_103) begin // @[ReservationStation.scala 83:7]
      if (reservation_2_valid) begin // @[ReservationStation.scala 85:27]
        reservation_2_ready1 <= _GEN_971;
      end else begin
        reservation_2_ready1 <= _GEN_931;
      end
    end else begin
      reservation_2_ready1 <= _GEN_931;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_2_value1 <= 64'h0; // @[ReservationStation.scala 28:28]
    end else if (_T_103) begin // @[ReservationStation.scala 83:7]
      if (reservation_2_valid) begin // @[ReservationStation.scala 85:27]
        if (~reservation_2_ready1 & _T_127) begin // @[ReservationStation.scala 86:79]
          reservation_2_value1 <= io_collectedOutput_1_outputs_bits_value; // @[ReservationStation.scala 87:26]
        end else begin
          reservation_2_value1 <= _GEN_930;
        end
      end else begin
        reservation_2_value1 <= _GEN_930;
      end
    end else begin
      reservation_2_value1 <= _GEN_930;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_2_sourceTag2_threadId <= 1'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h2 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_2_sourceTag2_threadId <= io_decoder_1_entry_sourceTag2_threadId; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_2_sourceTag2_threadId <= _GEN_427;
        end
      end else begin
        reservation_2_sourceTag2_threadId <= _GEN_427;
      end
    end else begin
      reservation_2_sourceTag2_threadId <= _GEN_427;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_2_sourceTag2_id <= 4'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h2 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_2_sourceTag2_id <= io_decoder_1_entry_sourceTag2_id; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_2_sourceTag2_id <= _GEN_435;
        end
      end else begin
        reservation_2_sourceTag2_id <= _GEN_435;
      end
    end else begin
      reservation_2_sourceTag2_id <= _GEN_435;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_2_ready2 <= 1'h0; // @[ReservationStation.scala 28:28]
    end else if (_T_103) begin // @[ReservationStation.scala 83:7]
      if (reservation_2_valid) begin // @[ReservationStation.scala 85:27]
        reservation_2_ready2 <= _GEN_973;
      end else begin
        reservation_2_ready2 <= _GEN_933;
      end
    end else begin
      reservation_2_ready2 <= _GEN_933;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_2_value2 <= 64'h0; // @[ReservationStation.scala 28:28]
    end else if (_T_103) begin // @[ReservationStation.scala 83:7]
      if (reservation_2_valid) begin // @[ReservationStation.scala 85:27]
        if (~reservation_2_ready2 & _T_132) begin // @[ReservationStation.scala 90:79]
          reservation_2_value2 <= io_collectedOutput_1_outputs_bits_value; // @[ReservationStation.scala 91:26]
        end else begin
          reservation_2_value2 <= _GEN_932;
        end
      end else begin
        reservation_2_value2 <= _GEN_932;
      end
    end else begin
      reservation_2_value2 <= _GEN_932;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_2_destinationTag_threadId <= 1'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        reservation_2_destinationTag_threadId <= _GEN_587;
      end else begin
        reservation_2_destinationTag_threadId <= _GEN_459;
      end
    end else begin
      reservation_2_destinationTag_threadId <= _GEN_459;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_2_destinationTag_id <= 4'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h2 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_2_destinationTag_id <= io_decoder_1_entry_destinationTag_id; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_2_destinationTag_id <= _GEN_467;
        end
      end else begin
        reservation_2_destinationTag_id <= _GEN_467;
      end
    end else begin
      reservation_2_destinationTag_id <= _GEN_467;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_2_wasCompressed <= 1'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h2 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_2_wasCompressed <= io_decoder_1_entry_wasCompressed; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_2_wasCompressed <= _GEN_475;
        end
      end else begin
        reservation_2_wasCompressed <= _GEN_475;
      end
    end else begin
      reservation_2_wasCompressed <= _GEN_475;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_2_valid <= 1'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h2 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_2_valid <= io_decoder_1_entry_valid; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_2_valid <= _GEN_483;
        end
      end else begin
        reservation_2_valid <= _GEN_483;
      end
    end else begin
      reservation_2_valid <= _GEN_483;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_3_opcode <= 7'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h3 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_3_opcode <= io_decoder_1_entry_opcode; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_3_opcode <= _GEN_372;
        end
      end else begin
        reservation_3_opcode <= _GEN_372;
      end
    end else begin
      reservation_3_opcode <= _GEN_372;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_3_function3 <= 3'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h3 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_3_function3 <= io_decoder_1_entry_function3; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_3_function3 <= _GEN_380;
        end
      end else begin
        reservation_3_function3 <= _GEN_380;
      end
    end else begin
      reservation_3_function3 <= _GEN_380;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_3_immediateOrFunction7 <= 12'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h3 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_3_immediateOrFunction7 <= io_decoder_1_entry_immediateOrFunction7; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_3_immediateOrFunction7 <= _GEN_388;
        end
      end else begin
        reservation_3_immediateOrFunction7 <= _GEN_388;
      end
    end else begin
      reservation_3_immediateOrFunction7 <= _GEN_388;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_3_sourceTag1_threadId <= 1'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h3 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_3_sourceTag1_threadId <= io_decoder_1_entry_sourceTag1_threadId; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_3_sourceTag1_threadId <= _GEN_396;
        end
      end else begin
        reservation_3_sourceTag1_threadId <= _GEN_396;
      end
    end else begin
      reservation_3_sourceTag1_threadId <= _GEN_396;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_3_sourceTag1_id <= 4'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h3 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_3_sourceTag1_id <= io_decoder_1_entry_sourceTag1_id; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_3_sourceTag1_id <= _GEN_404;
        end
      end else begin
        reservation_3_sourceTag1_id <= _GEN_404;
      end
    end else begin
      reservation_3_sourceTag1_id <= _GEN_404;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_3_ready1 <= 1'h0; // @[ReservationStation.scala 28:28]
    end else if (_T_103) begin // @[ReservationStation.scala 83:7]
      if (reservation_3_valid) begin // @[ReservationStation.scala 85:27]
        reservation_3_ready1 <= _GEN_979;
      end else begin
        reservation_3_ready1 <= _GEN_935;
      end
    end else begin
      reservation_3_ready1 <= _GEN_935;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_3_value1 <= 64'h0; // @[ReservationStation.scala 28:28]
    end else if (_T_103) begin // @[ReservationStation.scala 83:7]
      if (reservation_3_valid) begin // @[ReservationStation.scala 85:27]
        if (~reservation_3_ready1 & _T_137) begin // @[ReservationStation.scala 86:79]
          reservation_3_value1 <= io_collectedOutput_1_outputs_bits_value; // @[ReservationStation.scala 87:26]
        end else begin
          reservation_3_value1 <= _GEN_934;
        end
      end else begin
        reservation_3_value1 <= _GEN_934;
      end
    end else begin
      reservation_3_value1 <= _GEN_934;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_3_sourceTag2_threadId <= 1'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h3 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_3_sourceTag2_threadId <= io_decoder_1_entry_sourceTag2_threadId; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_3_sourceTag2_threadId <= _GEN_428;
        end
      end else begin
        reservation_3_sourceTag2_threadId <= _GEN_428;
      end
    end else begin
      reservation_3_sourceTag2_threadId <= _GEN_428;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_3_sourceTag2_id <= 4'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h3 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_3_sourceTag2_id <= io_decoder_1_entry_sourceTag2_id; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_3_sourceTag2_id <= _GEN_436;
        end
      end else begin
        reservation_3_sourceTag2_id <= _GEN_436;
      end
    end else begin
      reservation_3_sourceTag2_id <= _GEN_436;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_3_ready2 <= 1'h0; // @[ReservationStation.scala 28:28]
    end else if (_T_103) begin // @[ReservationStation.scala 83:7]
      if (reservation_3_valid) begin // @[ReservationStation.scala 85:27]
        reservation_3_ready2 <= _GEN_981;
      end else begin
        reservation_3_ready2 <= _GEN_937;
      end
    end else begin
      reservation_3_ready2 <= _GEN_937;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_3_value2 <= 64'h0; // @[ReservationStation.scala 28:28]
    end else if (_T_103) begin // @[ReservationStation.scala 83:7]
      if (reservation_3_valid) begin // @[ReservationStation.scala 85:27]
        if (~reservation_3_ready2 & _T_142) begin // @[ReservationStation.scala 90:79]
          reservation_3_value2 <= io_collectedOutput_1_outputs_bits_value; // @[ReservationStation.scala 91:26]
        end else begin
          reservation_3_value2 <= _GEN_936;
        end
      end else begin
        reservation_3_value2 <= _GEN_936;
      end
    end else begin
      reservation_3_value2 <= _GEN_936;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_3_destinationTag_threadId <= 1'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        reservation_3_destinationTag_threadId <= _GEN_588;
      end else begin
        reservation_3_destinationTag_threadId <= _GEN_460;
      end
    end else begin
      reservation_3_destinationTag_threadId <= _GEN_460;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_3_destinationTag_id <= 4'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h3 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_3_destinationTag_id <= io_decoder_1_entry_destinationTag_id; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_3_destinationTag_id <= _GEN_468;
        end
      end else begin
        reservation_3_destinationTag_id <= _GEN_468;
      end
    end else begin
      reservation_3_destinationTag_id <= _GEN_468;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_3_wasCompressed <= 1'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h3 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_3_wasCompressed <= io_decoder_1_entry_wasCompressed; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_3_wasCompressed <= _GEN_476;
        end
      end else begin
        reservation_3_wasCompressed <= _GEN_476;
      end
    end else begin
      reservation_3_wasCompressed <= _GEN_476;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_3_valid <= 1'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h3 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_3_valid <= io_decoder_1_entry_valid; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_3_valid <= _GEN_484;
        end
      end else begin
        reservation_3_valid <= _GEN_484;
      end
    end else begin
      reservation_3_valid <= _GEN_484;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_4_opcode <= 7'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h4 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_4_opcode <= io_decoder_1_entry_opcode; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_4_opcode <= _GEN_373;
        end
      end else begin
        reservation_4_opcode <= _GEN_373;
      end
    end else begin
      reservation_4_opcode <= _GEN_373;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_4_function3 <= 3'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h4 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_4_function3 <= io_decoder_1_entry_function3; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_4_function3 <= _GEN_381;
        end
      end else begin
        reservation_4_function3 <= _GEN_381;
      end
    end else begin
      reservation_4_function3 <= _GEN_381;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_4_immediateOrFunction7 <= 12'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h4 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_4_immediateOrFunction7 <= io_decoder_1_entry_immediateOrFunction7; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_4_immediateOrFunction7 <= _GEN_389;
        end
      end else begin
        reservation_4_immediateOrFunction7 <= _GEN_389;
      end
    end else begin
      reservation_4_immediateOrFunction7 <= _GEN_389;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_4_sourceTag1_threadId <= 1'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h4 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_4_sourceTag1_threadId <= io_decoder_1_entry_sourceTag1_threadId; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_4_sourceTag1_threadId <= _GEN_397;
        end
      end else begin
        reservation_4_sourceTag1_threadId <= _GEN_397;
      end
    end else begin
      reservation_4_sourceTag1_threadId <= _GEN_397;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_4_sourceTag1_id <= 4'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h4 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_4_sourceTag1_id <= io_decoder_1_entry_sourceTag1_id; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_4_sourceTag1_id <= _GEN_405;
        end
      end else begin
        reservation_4_sourceTag1_id <= _GEN_405;
      end
    end else begin
      reservation_4_sourceTag1_id <= _GEN_405;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_4_ready1 <= 1'h0; // @[ReservationStation.scala 28:28]
    end else if (_T_103) begin // @[ReservationStation.scala 83:7]
      if (reservation_4_valid) begin // @[ReservationStation.scala 85:27]
        reservation_4_ready1 <= _GEN_987;
      end else begin
        reservation_4_ready1 <= _GEN_939;
      end
    end else begin
      reservation_4_ready1 <= _GEN_939;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_4_value1 <= 64'h0; // @[ReservationStation.scala 28:28]
    end else if (_T_103) begin // @[ReservationStation.scala 83:7]
      if (reservation_4_valid) begin // @[ReservationStation.scala 85:27]
        if (~reservation_4_ready1 & _T_147) begin // @[ReservationStation.scala 86:79]
          reservation_4_value1 <= io_collectedOutput_1_outputs_bits_value; // @[ReservationStation.scala 87:26]
        end else begin
          reservation_4_value1 <= _GEN_938;
        end
      end else begin
        reservation_4_value1 <= _GEN_938;
      end
    end else begin
      reservation_4_value1 <= _GEN_938;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_4_sourceTag2_threadId <= 1'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h4 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_4_sourceTag2_threadId <= io_decoder_1_entry_sourceTag2_threadId; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_4_sourceTag2_threadId <= _GEN_429;
        end
      end else begin
        reservation_4_sourceTag2_threadId <= _GEN_429;
      end
    end else begin
      reservation_4_sourceTag2_threadId <= _GEN_429;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_4_sourceTag2_id <= 4'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h4 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_4_sourceTag2_id <= io_decoder_1_entry_sourceTag2_id; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_4_sourceTag2_id <= _GEN_437;
        end
      end else begin
        reservation_4_sourceTag2_id <= _GEN_437;
      end
    end else begin
      reservation_4_sourceTag2_id <= _GEN_437;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_4_ready2 <= 1'h0; // @[ReservationStation.scala 28:28]
    end else if (_T_103) begin // @[ReservationStation.scala 83:7]
      if (reservation_4_valid) begin // @[ReservationStation.scala 85:27]
        reservation_4_ready2 <= _GEN_989;
      end else begin
        reservation_4_ready2 <= _GEN_941;
      end
    end else begin
      reservation_4_ready2 <= _GEN_941;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_4_value2 <= 64'h0; // @[ReservationStation.scala 28:28]
    end else if (_T_103) begin // @[ReservationStation.scala 83:7]
      if (reservation_4_valid) begin // @[ReservationStation.scala 85:27]
        if (~reservation_4_ready2 & _T_152) begin // @[ReservationStation.scala 90:79]
          reservation_4_value2 <= io_collectedOutput_1_outputs_bits_value; // @[ReservationStation.scala 91:26]
        end else begin
          reservation_4_value2 <= _GEN_940;
        end
      end else begin
        reservation_4_value2 <= _GEN_940;
      end
    end else begin
      reservation_4_value2 <= _GEN_940;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_4_destinationTag_threadId <= 1'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        reservation_4_destinationTag_threadId <= _GEN_589;
      end else begin
        reservation_4_destinationTag_threadId <= _GEN_461;
      end
    end else begin
      reservation_4_destinationTag_threadId <= _GEN_461;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_4_destinationTag_id <= 4'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h4 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_4_destinationTag_id <= io_decoder_1_entry_destinationTag_id; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_4_destinationTag_id <= _GEN_469;
        end
      end else begin
        reservation_4_destinationTag_id <= _GEN_469;
      end
    end else begin
      reservation_4_destinationTag_id <= _GEN_469;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_4_wasCompressed <= 1'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h4 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_4_wasCompressed <= io_decoder_1_entry_wasCompressed; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_4_wasCompressed <= _GEN_477;
        end
      end else begin
        reservation_4_wasCompressed <= _GEN_477;
      end
    end else begin
      reservation_4_wasCompressed <= _GEN_477;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_4_valid <= 1'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h4 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_4_valid <= io_decoder_1_entry_valid; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_4_valid <= _GEN_485;
        end
      end else begin
        reservation_4_valid <= _GEN_485;
      end
    end else begin
      reservation_4_valid <= _GEN_485;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_5_opcode <= 7'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h5 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_5_opcode <= io_decoder_1_entry_opcode; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_5_opcode <= _GEN_374;
        end
      end else begin
        reservation_5_opcode <= _GEN_374;
      end
    end else begin
      reservation_5_opcode <= _GEN_374;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_5_function3 <= 3'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h5 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_5_function3 <= io_decoder_1_entry_function3; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_5_function3 <= _GEN_382;
        end
      end else begin
        reservation_5_function3 <= _GEN_382;
      end
    end else begin
      reservation_5_function3 <= _GEN_382;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_5_immediateOrFunction7 <= 12'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h5 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_5_immediateOrFunction7 <= io_decoder_1_entry_immediateOrFunction7; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_5_immediateOrFunction7 <= _GEN_390;
        end
      end else begin
        reservation_5_immediateOrFunction7 <= _GEN_390;
      end
    end else begin
      reservation_5_immediateOrFunction7 <= _GEN_390;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_5_sourceTag1_threadId <= 1'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h5 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_5_sourceTag1_threadId <= io_decoder_1_entry_sourceTag1_threadId; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_5_sourceTag1_threadId <= _GEN_398;
        end
      end else begin
        reservation_5_sourceTag1_threadId <= _GEN_398;
      end
    end else begin
      reservation_5_sourceTag1_threadId <= _GEN_398;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_5_sourceTag1_id <= 4'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h5 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_5_sourceTag1_id <= io_decoder_1_entry_sourceTag1_id; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_5_sourceTag1_id <= _GEN_406;
        end
      end else begin
        reservation_5_sourceTag1_id <= _GEN_406;
      end
    end else begin
      reservation_5_sourceTag1_id <= _GEN_406;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_5_ready1 <= 1'h0; // @[ReservationStation.scala 28:28]
    end else if (_T_103) begin // @[ReservationStation.scala 83:7]
      if (reservation_5_valid) begin // @[ReservationStation.scala 85:27]
        reservation_5_ready1 <= _GEN_995;
      end else begin
        reservation_5_ready1 <= _GEN_943;
      end
    end else begin
      reservation_5_ready1 <= _GEN_943;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_5_value1 <= 64'h0; // @[ReservationStation.scala 28:28]
    end else if (_T_103) begin // @[ReservationStation.scala 83:7]
      if (reservation_5_valid) begin // @[ReservationStation.scala 85:27]
        if (~reservation_5_ready1 & _T_157) begin // @[ReservationStation.scala 86:79]
          reservation_5_value1 <= io_collectedOutput_1_outputs_bits_value; // @[ReservationStation.scala 87:26]
        end else begin
          reservation_5_value1 <= _GEN_942;
        end
      end else begin
        reservation_5_value1 <= _GEN_942;
      end
    end else begin
      reservation_5_value1 <= _GEN_942;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_5_sourceTag2_threadId <= 1'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h5 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_5_sourceTag2_threadId <= io_decoder_1_entry_sourceTag2_threadId; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_5_sourceTag2_threadId <= _GEN_430;
        end
      end else begin
        reservation_5_sourceTag2_threadId <= _GEN_430;
      end
    end else begin
      reservation_5_sourceTag2_threadId <= _GEN_430;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_5_sourceTag2_id <= 4'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h5 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_5_sourceTag2_id <= io_decoder_1_entry_sourceTag2_id; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_5_sourceTag2_id <= _GEN_438;
        end
      end else begin
        reservation_5_sourceTag2_id <= _GEN_438;
      end
    end else begin
      reservation_5_sourceTag2_id <= _GEN_438;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_5_ready2 <= 1'h0; // @[ReservationStation.scala 28:28]
    end else if (_T_103) begin // @[ReservationStation.scala 83:7]
      if (reservation_5_valid) begin // @[ReservationStation.scala 85:27]
        reservation_5_ready2 <= _GEN_997;
      end else begin
        reservation_5_ready2 <= _GEN_945;
      end
    end else begin
      reservation_5_ready2 <= _GEN_945;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_5_value2 <= 64'h0; // @[ReservationStation.scala 28:28]
    end else if (_T_103) begin // @[ReservationStation.scala 83:7]
      if (reservation_5_valid) begin // @[ReservationStation.scala 85:27]
        if (~reservation_5_ready2 & _T_162) begin // @[ReservationStation.scala 90:79]
          reservation_5_value2 <= io_collectedOutput_1_outputs_bits_value; // @[ReservationStation.scala 91:26]
        end else begin
          reservation_5_value2 <= _GEN_944;
        end
      end else begin
        reservation_5_value2 <= _GEN_944;
      end
    end else begin
      reservation_5_value2 <= _GEN_944;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_5_destinationTag_threadId <= 1'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        reservation_5_destinationTag_threadId <= _GEN_590;
      end else begin
        reservation_5_destinationTag_threadId <= _GEN_462;
      end
    end else begin
      reservation_5_destinationTag_threadId <= _GEN_462;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_5_destinationTag_id <= 4'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h5 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_5_destinationTag_id <= io_decoder_1_entry_destinationTag_id; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_5_destinationTag_id <= _GEN_470;
        end
      end else begin
        reservation_5_destinationTag_id <= _GEN_470;
      end
    end else begin
      reservation_5_destinationTag_id <= _GEN_470;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_5_wasCompressed <= 1'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h5 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_5_wasCompressed <= io_decoder_1_entry_wasCompressed; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_5_wasCompressed <= _GEN_478;
        end
      end else begin
        reservation_5_wasCompressed <= _GEN_478;
      end
    end else begin
      reservation_5_wasCompressed <= _GEN_478;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_5_valid <= 1'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h5 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_5_valid <= io_decoder_1_entry_valid; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_5_valid <= _GEN_486;
        end
      end else begin
        reservation_5_valid <= _GEN_486;
      end
    end else begin
      reservation_5_valid <= _GEN_486;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_6_opcode <= 7'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h6 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_6_opcode <= io_decoder_1_entry_opcode; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_6_opcode <= _GEN_375;
        end
      end else begin
        reservation_6_opcode <= _GEN_375;
      end
    end else begin
      reservation_6_opcode <= _GEN_375;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_6_function3 <= 3'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h6 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_6_function3 <= io_decoder_1_entry_function3; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_6_function3 <= _GEN_383;
        end
      end else begin
        reservation_6_function3 <= _GEN_383;
      end
    end else begin
      reservation_6_function3 <= _GEN_383;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_6_immediateOrFunction7 <= 12'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h6 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_6_immediateOrFunction7 <= io_decoder_1_entry_immediateOrFunction7; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_6_immediateOrFunction7 <= _GEN_391;
        end
      end else begin
        reservation_6_immediateOrFunction7 <= _GEN_391;
      end
    end else begin
      reservation_6_immediateOrFunction7 <= _GEN_391;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_6_sourceTag1_threadId <= 1'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h6 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_6_sourceTag1_threadId <= io_decoder_1_entry_sourceTag1_threadId; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_6_sourceTag1_threadId <= _GEN_399;
        end
      end else begin
        reservation_6_sourceTag1_threadId <= _GEN_399;
      end
    end else begin
      reservation_6_sourceTag1_threadId <= _GEN_399;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_6_sourceTag1_id <= 4'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h6 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_6_sourceTag1_id <= io_decoder_1_entry_sourceTag1_id; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_6_sourceTag1_id <= _GEN_407;
        end
      end else begin
        reservation_6_sourceTag1_id <= _GEN_407;
      end
    end else begin
      reservation_6_sourceTag1_id <= _GEN_407;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_6_ready1 <= 1'h0; // @[ReservationStation.scala 28:28]
    end else if (_T_103) begin // @[ReservationStation.scala 83:7]
      if (reservation_6_valid) begin // @[ReservationStation.scala 85:27]
        reservation_6_ready1 <= _GEN_1003;
      end else begin
        reservation_6_ready1 <= _GEN_947;
      end
    end else begin
      reservation_6_ready1 <= _GEN_947;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_6_value1 <= 64'h0; // @[ReservationStation.scala 28:28]
    end else if (_T_103) begin // @[ReservationStation.scala 83:7]
      if (reservation_6_valid) begin // @[ReservationStation.scala 85:27]
        if (~reservation_6_ready1 & _T_167) begin // @[ReservationStation.scala 86:79]
          reservation_6_value1 <= io_collectedOutput_1_outputs_bits_value; // @[ReservationStation.scala 87:26]
        end else begin
          reservation_6_value1 <= _GEN_946;
        end
      end else begin
        reservation_6_value1 <= _GEN_946;
      end
    end else begin
      reservation_6_value1 <= _GEN_946;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_6_sourceTag2_threadId <= 1'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h6 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_6_sourceTag2_threadId <= io_decoder_1_entry_sourceTag2_threadId; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_6_sourceTag2_threadId <= _GEN_431;
        end
      end else begin
        reservation_6_sourceTag2_threadId <= _GEN_431;
      end
    end else begin
      reservation_6_sourceTag2_threadId <= _GEN_431;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_6_sourceTag2_id <= 4'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h6 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_6_sourceTag2_id <= io_decoder_1_entry_sourceTag2_id; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_6_sourceTag2_id <= _GEN_439;
        end
      end else begin
        reservation_6_sourceTag2_id <= _GEN_439;
      end
    end else begin
      reservation_6_sourceTag2_id <= _GEN_439;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_6_ready2 <= 1'h0; // @[ReservationStation.scala 28:28]
    end else if (_T_103) begin // @[ReservationStation.scala 83:7]
      if (reservation_6_valid) begin // @[ReservationStation.scala 85:27]
        reservation_6_ready2 <= _GEN_1005;
      end else begin
        reservation_6_ready2 <= _GEN_949;
      end
    end else begin
      reservation_6_ready2 <= _GEN_949;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_6_value2 <= 64'h0; // @[ReservationStation.scala 28:28]
    end else if (_T_103) begin // @[ReservationStation.scala 83:7]
      if (reservation_6_valid) begin // @[ReservationStation.scala 85:27]
        if (~reservation_6_ready2 & _T_172) begin // @[ReservationStation.scala 90:79]
          reservation_6_value2 <= io_collectedOutput_1_outputs_bits_value; // @[ReservationStation.scala 91:26]
        end else begin
          reservation_6_value2 <= _GEN_948;
        end
      end else begin
        reservation_6_value2 <= _GEN_948;
      end
    end else begin
      reservation_6_value2 <= _GEN_948;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_6_destinationTag_threadId <= 1'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        reservation_6_destinationTag_threadId <= _GEN_591;
      end else begin
        reservation_6_destinationTag_threadId <= _GEN_463;
      end
    end else begin
      reservation_6_destinationTag_threadId <= _GEN_463;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_6_destinationTag_id <= 4'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h6 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_6_destinationTag_id <= io_decoder_1_entry_destinationTag_id; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_6_destinationTag_id <= _GEN_471;
        end
      end else begin
        reservation_6_destinationTag_id <= _GEN_471;
      end
    end else begin
      reservation_6_destinationTag_id <= _GEN_471;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_6_wasCompressed <= 1'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h6 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_6_wasCompressed <= io_decoder_1_entry_wasCompressed; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_6_wasCompressed <= _GEN_479;
        end
      end else begin
        reservation_6_wasCompressed <= _GEN_479;
      end
    end else begin
      reservation_6_wasCompressed <= _GEN_479;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_6_valid <= 1'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h6 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_6_valid <= io_decoder_1_entry_valid; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_6_valid <= _GEN_487;
        end
      end else begin
        reservation_6_valid <= _GEN_487;
      end
    end else begin
      reservation_6_valid <= _GEN_487;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_7_opcode <= 7'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h7 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_7_opcode <= io_decoder_1_entry_opcode; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_7_opcode <= _GEN_376;
        end
      end else begin
        reservation_7_opcode <= _GEN_376;
      end
    end else begin
      reservation_7_opcode <= _GEN_376;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_7_function3 <= 3'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h7 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_7_function3 <= io_decoder_1_entry_function3; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_7_function3 <= _GEN_384;
        end
      end else begin
        reservation_7_function3 <= _GEN_384;
      end
    end else begin
      reservation_7_function3 <= _GEN_384;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_7_immediateOrFunction7 <= 12'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h7 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_7_immediateOrFunction7 <= io_decoder_1_entry_immediateOrFunction7; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_7_immediateOrFunction7 <= _GEN_392;
        end
      end else begin
        reservation_7_immediateOrFunction7 <= _GEN_392;
      end
    end else begin
      reservation_7_immediateOrFunction7 <= _GEN_392;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_7_sourceTag1_threadId <= 1'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h7 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_7_sourceTag1_threadId <= io_decoder_1_entry_sourceTag1_threadId; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_7_sourceTag1_threadId <= _GEN_400;
        end
      end else begin
        reservation_7_sourceTag1_threadId <= _GEN_400;
      end
    end else begin
      reservation_7_sourceTag1_threadId <= _GEN_400;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_7_sourceTag1_id <= 4'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h7 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_7_sourceTag1_id <= io_decoder_1_entry_sourceTag1_id; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_7_sourceTag1_id <= _GEN_408;
        end
      end else begin
        reservation_7_sourceTag1_id <= _GEN_408;
      end
    end else begin
      reservation_7_sourceTag1_id <= _GEN_408;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_7_ready1 <= 1'h0; // @[ReservationStation.scala 28:28]
    end else if (_T_103) begin // @[ReservationStation.scala 83:7]
      if (reservation_7_valid) begin // @[ReservationStation.scala 85:27]
        reservation_7_ready1 <= _GEN_1011;
      end else begin
        reservation_7_ready1 <= _GEN_951;
      end
    end else begin
      reservation_7_ready1 <= _GEN_951;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_7_value1 <= 64'h0; // @[ReservationStation.scala 28:28]
    end else if (_T_103) begin // @[ReservationStation.scala 83:7]
      if (reservation_7_valid) begin // @[ReservationStation.scala 85:27]
        if (~reservation_7_ready1 & _T_177) begin // @[ReservationStation.scala 86:79]
          reservation_7_value1 <= io_collectedOutput_1_outputs_bits_value; // @[ReservationStation.scala 87:26]
        end else begin
          reservation_7_value1 <= _GEN_950;
        end
      end else begin
        reservation_7_value1 <= _GEN_950;
      end
    end else begin
      reservation_7_value1 <= _GEN_950;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_7_sourceTag2_threadId <= 1'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h7 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_7_sourceTag2_threadId <= io_decoder_1_entry_sourceTag2_threadId; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_7_sourceTag2_threadId <= _GEN_432;
        end
      end else begin
        reservation_7_sourceTag2_threadId <= _GEN_432;
      end
    end else begin
      reservation_7_sourceTag2_threadId <= _GEN_432;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_7_sourceTag2_id <= 4'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h7 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_7_sourceTag2_id <= io_decoder_1_entry_sourceTag2_id; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_7_sourceTag2_id <= _GEN_440;
        end
      end else begin
        reservation_7_sourceTag2_id <= _GEN_440;
      end
    end else begin
      reservation_7_sourceTag2_id <= _GEN_440;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_7_ready2 <= 1'h0; // @[ReservationStation.scala 28:28]
    end else if (_T_103) begin // @[ReservationStation.scala 83:7]
      if (reservation_7_valid) begin // @[ReservationStation.scala 85:27]
        reservation_7_ready2 <= _GEN_1013;
      end else begin
        reservation_7_ready2 <= _GEN_953;
      end
    end else begin
      reservation_7_ready2 <= _GEN_953;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_7_value2 <= 64'h0; // @[ReservationStation.scala 28:28]
    end else if (_T_103) begin // @[ReservationStation.scala 83:7]
      if (reservation_7_valid) begin // @[ReservationStation.scala 85:27]
        if (~reservation_7_ready2 & _T_182) begin // @[ReservationStation.scala 90:79]
          reservation_7_value2 <= io_collectedOutput_1_outputs_bits_value; // @[ReservationStation.scala 91:26]
        end else begin
          reservation_7_value2 <= _GEN_952;
        end
      end else begin
        reservation_7_value2 <= _GEN_952;
      end
    end else begin
      reservation_7_value2 <= _GEN_952;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_7_destinationTag_threadId <= 1'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        reservation_7_destinationTag_threadId <= _GEN_592;
      end else begin
        reservation_7_destinationTag_threadId <= _GEN_464;
      end
    end else begin
      reservation_7_destinationTag_threadId <= _GEN_464;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_7_destinationTag_id <= 4'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h7 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_7_destinationTag_id <= io_decoder_1_entry_destinationTag_id; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_7_destinationTag_id <= _GEN_472;
        end
      end else begin
        reservation_7_destinationTag_id <= _GEN_472;
      end
    end else begin
      reservation_7_destinationTag_id <= _GEN_472;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_7_wasCompressed <= 1'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h7 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_7_wasCompressed <= io_decoder_1_entry_wasCompressed; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_7_wasCompressed <= _GEN_480;
        end
      end else begin
        reservation_7_wasCompressed <= _GEN_480;
      end
    end else begin
      reservation_7_wasCompressed <= _GEN_480;
    end
    if (reset) begin // @[ReservationStation.scala 28:28]
      reservation_7_valid <= 1'h0; // @[ReservationStation.scala 28:28]
    end else if (~_GEN_496) begin // @[ReservationStation.scala 66:40]
      if (io_decoder_1_entry_valid) begin // @[ReservationStation.scala 68:39]
        if (3'h7 == _T_13) begin // @[ReservationStation.scala 69:31]
          reservation_7_valid <= io_decoder_1_entry_valid; // @[ReservationStation.scala 69:31]
        end else begin
          reservation_7_valid <= _GEN_488;
        end
      end else begin
        reservation_7_valid <= _GEN_488;
      end
    end else begin
      reservation_7_valid <= _GEN_488;
    end
    if (reset) begin // @[ReservationStation.scala 62:29]
      head <= 3'h0; // @[ReservationStation.scala 62:29]
    end else if (_T_16) begin // @[ReservationStation.scala 72:19]
      head <= _T_18;
    end else if (_T_10) begin // @[ReservationStation.scala 72:19]
      head <= _T_12;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reservation_0_opcode = _RAND_0[6:0];
  _RAND_1 = {1{`RANDOM}};
  reservation_0_function3 = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  reservation_0_immediateOrFunction7 = _RAND_2[11:0];
  _RAND_3 = {1{`RANDOM}};
  reservation_0_sourceTag1_threadId = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  reservation_0_sourceTag1_id = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  reservation_0_ready1 = _RAND_5[0:0];
  _RAND_6 = {2{`RANDOM}};
  reservation_0_value1 = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  reservation_0_sourceTag2_threadId = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  reservation_0_sourceTag2_id = _RAND_8[3:0];
  _RAND_9 = {1{`RANDOM}};
  reservation_0_ready2 = _RAND_9[0:0];
  _RAND_10 = {2{`RANDOM}};
  reservation_0_value2 = _RAND_10[63:0];
  _RAND_11 = {1{`RANDOM}};
  reservation_0_destinationTag_threadId = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  reservation_0_destinationTag_id = _RAND_12[3:0];
  _RAND_13 = {1{`RANDOM}};
  reservation_0_wasCompressed = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  reservation_0_valid = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  reservation_1_opcode = _RAND_15[6:0];
  _RAND_16 = {1{`RANDOM}};
  reservation_1_function3 = _RAND_16[2:0];
  _RAND_17 = {1{`RANDOM}};
  reservation_1_immediateOrFunction7 = _RAND_17[11:0];
  _RAND_18 = {1{`RANDOM}};
  reservation_1_sourceTag1_threadId = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  reservation_1_sourceTag1_id = _RAND_19[3:0];
  _RAND_20 = {1{`RANDOM}};
  reservation_1_ready1 = _RAND_20[0:0];
  _RAND_21 = {2{`RANDOM}};
  reservation_1_value1 = _RAND_21[63:0];
  _RAND_22 = {1{`RANDOM}};
  reservation_1_sourceTag2_threadId = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  reservation_1_sourceTag2_id = _RAND_23[3:0];
  _RAND_24 = {1{`RANDOM}};
  reservation_1_ready2 = _RAND_24[0:0];
  _RAND_25 = {2{`RANDOM}};
  reservation_1_value2 = _RAND_25[63:0];
  _RAND_26 = {1{`RANDOM}};
  reservation_1_destinationTag_threadId = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  reservation_1_destinationTag_id = _RAND_27[3:0];
  _RAND_28 = {1{`RANDOM}};
  reservation_1_wasCompressed = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  reservation_1_valid = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  reservation_2_opcode = _RAND_30[6:0];
  _RAND_31 = {1{`RANDOM}};
  reservation_2_function3 = _RAND_31[2:0];
  _RAND_32 = {1{`RANDOM}};
  reservation_2_immediateOrFunction7 = _RAND_32[11:0];
  _RAND_33 = {1{`RANDOM}};
  reservation_2_sourceTag1_threadId = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  reservation_2_sourceTag1_id = _RAND_34[3:0];
  _RAND_35 = {1{`RANDOM}};
  reservation_2_ready1 = _RAND_35[0:0];
  _RAND_36 = {2{`RANDOM}};
  reservation_2_value1 = _RAND_36[63:0];
  _RAND_37 = {1{`RANDOM}};
  reservation_2_sourceTag2_threadId = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  reservation_2_sourceTag2_id = _RAND_38[3:0];
  _RAND_39 = {1{`RANDOM}};
  reservation_2_ready2 = _RAND_39[0:0];
  _RAND_40 = {2{`RANDOM}};
  reservation_2_value2 = _RAND_40[63:0];
  _RAND_41 = {1{`RANDOM}};
  reservation_2_destinationTag_threadId = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  reservation_2_destinationTag_id = _RAND_42[3:0];
  _RAND_43 = {1{`RANDOM}};
  reservation_2_wasCompressed = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  reservation_2_valid = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  reservation_3_opcode = _RAND_45[6:0];
  _RAND_46 = {1{`RANDOM}};
  reservation_3_function3 = _RAND_46[2:0];
  _RAND_47 = {1{`RANDOM}};
  reservation_3_immediateOrFunction7 = _RAND_47[11:0];
  _RAND_48 = {1{`RANDOM}};
  reservation_3_sourceTag1_threadId = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  reservation_3_sourceTag1_id = _RAND_49[3:0];
  _RAND_50 = {1{`RANDOM}};
  reservation_3_ready1 = _RAND_50[0:0];
  _RAND_51 = {2{`RANDOM}};
  reservation_3_value1 = _RAND_51[63:0];
  _RAND_52 = {1{`RANDOM}};
  reservation_3_sourceTag2_threadId = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  reservation_3_sourceTag2_id = _RAND_53[3:0];
  _RAND_54 = {1{`RANDOM}};
  reservation_3_ready2 = _RAND_54[0:0];
  _RAND_55 = {2{`RANDOM}};
  reservation_3_value2 = _RAND_55[63:0];
  _RAND_56 = {1{`RANDOM}};
  reservation_3_destinationTag_threadId = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  reservation_3_destinationTag_id = _RAND_57[3:0];
  _RAND_58 = {1{`RANDOM}};
  reservation_3_wasCompressed = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  reservation_3_valid = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  reservation_4_opcode = _RAND_60[6:0];
  _RAND_61 = {1{`RANDOM}};
  reservation_4_function3 = _RAND_61[2:0];
  _RAND_62 = {1{`RANDOM}};
  reservation_4_immediateOrFunction7 = _RAND_62[11:0];
  _RAND_63 = {1{`RANDOM}};
  reservation_4_sourceTag1_threadId = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  reservation_4_sourceTag1_id = _RAND_64[3:0];
  _RAND_65 = {1{`RANDOM}};
  reservation_4_ready1 = _RAND_65[0:0];
  _RAND_66 = {2{`RANDOM}};
  reservation_4_value1 = _RAND_66[63:0];
  _RAND_67 = {1{`RANDOM}};
  reservation_4_sourceTag2_threadId = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  reservation_4_sourceTag2_id = _RAND_68[3:0];
  _RAND_69 = {1{`RANDOM}};
  reservation_4_ready2 = _RAND_69[0:0];
  _RAND_70 = {2{`RANDOM}};
  reservation_4_value2 = _RAND_70[63:0];
  _RAND_71 = {1{`RANDOM}};
  reservation_4_destinationTag_threadId = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  reservation_4_destinationTag_id = _RAND_72[3:0];
  _RAND_73 = {1{`RANDOM}};
  reservation_4_wasCompressed = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  reservation_4_valid = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  reservation_5_opcode = _RAND_75[6:0];
  _RAND_76 = {1{`RANDOM}};
  reservation_5_function3 = _RAND_76[2:0];
  _RAND_77 = {1{`RANDOM}};
  reservation_5_immediateOrFunction7 = _RAND_77[11:0];
  _RAND_78 = {1{`RANDOM}};
  reservation_5_sourceTag1_threadId = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  reservation_5_sourceTag1_id = _RAND_79[3:0];
  _RAND_80 = {1{`RANDOM}};
  reservation_5_ready1 = _RAND_80[0:0];
  _RAND_81 = {2{`RANDOM}};
  reservation_5_value1 = _RAND_81[63:0];
  _RAND_82 = {1{`RANDOM}};
  reservation_5_sourceTag2_threadId = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  reservation_5_sourceTag2_id = _RAND_83[3:0];
  _RAND_84 = {1{`RANDOM}};
  reservation_5_ready2 = _RAND_84[0:0];
  _RAND_85 = {2{`RANDOM}};
  reservation_5_value2 = _RAND_85[63:0];
  _RAND_86 = {1{`RANDOM}};
  reservation_5_destinationTag_threadId = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  reservation_5_destinationTag_id = _RAND_87[3:0];
  _RAND_88 = {1{`RANDOM}};
  reservation_5_wasCompressed = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  reservation_5_valid = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  reservation_6_opcode = _RAND_90[6:0];
  _RAND_91 = {1{`RANDOM}};
  reservation_6_function3 = _RAND_91[2:0];
  _RAND_92 = {1{`RANDOM}};
  reservation_6_immediateOrFunction7 = _RAND_92[11:0];
  _RAND_93 = {1{`RANDOM}};
  reservation_6_sourceTag1_threadId = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  reservation_6_sourceTag1_id = _RAND_94[3:0];
  _RAND_95 = {1{`RANDOM}};
  reservation_6_ready1 = _RAND_95[0:0];
  _RAND_96 = {2{`RANDOM}};
  reservation_6_value1 = _RAND_96[63:0];
  _RAND_97 = {1{`RANDOM}};
  reservation_6_sourceTag2_threadId = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  reservation_6_sourceTag2_id = _RAND_98[3:0];
  _RAND_99 = {1{`RANDOM}};
  reservation_6_ready2 = _RAND_99[0:0];
  _RAND_100 = {2{`RANDOM}};
  reservation_6_value2 = _RAND_100[63:0];
  _RAND_101 = {1{`RANDOM}};
  reservation_6_destinationTag_threadId = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  reservation_6_destinationTag_id = _RAND_102[3:0];
  _RAND_103 = {1{`RANDOM}};
  reservation_6_wasCompressed = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  reservation_6_valid = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  reservation_7_opcode = _RAND_105[6:0];
  _RAND_106 = {1{`RANDOM}};
  reservation_7_function3 = _RAND_106[2:0];
  _RAND_107 = {1{`RANDOM}};
  reservation_7_immediateOrFunction7 = _RAND_107[11:0];
  _RAND_108 = {1{`RANDOM}};
  reservation_7_sourceTag1_threadId = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  reservation_7_sourceTag1_id = _RAND_109[3:0];
  _RAND_110 = {1{`RANDOM}};
  reservation_7_ready1 = _RAND_110[0:0];
  _RAND_111 = {2{`RANDOM}};
  reservation_7_value1 = _RAND_111[63:0];
  _RAND_112 = {1{`RANDOM}};
  reservation_7_sourceTag2_threadId = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  reservation_7_sourceTag2_id = _RAND_113[3:0];
  _RAND_114 = {1{`RANDOM}};
  reservation_7_ready2 = _RAND_114[0:0];
  _RAND_115 = {2{`RANDOM}};
  reservation_7_value2 = _RAND_115[63:0];
  _RAND_116 = {1{`RANDOM}};
  reservation_7_destinationTag_threadId = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  reservation_7_destinationTag_id = _RAND_117[3:0];
  _RAND_118 = {1{`RANDOM}};
  reservation_7_wasCompressed = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  reservation_7_valid = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  head = _RAND_120[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module InstructionChecker(
  input  [2:0] input_function3bits,
  input  [6:0] input_function7bits,
  input  [6:0] input_opcode,
  output [3:0] output_instruction,
  output [2:0] output_branch,
  output [2:0] output_operationWidth,
  output [3:0] output_arithmetic
);
  wire [3:0] _output_instruction_T_1 = input_function3bits[0] ? 4'ha : 4'h9; // @[InstructionChecker.scala 27:26]
  wire  _output_instruction_T_2 = |input_function3bits; // @[InstructionChecker.scala 33:29]
  wire [3:0] _output_instruction_T_4 = input_function3bits[2] ? 4'he : 4'hd; // @[InstructionChecker.scala 34:12]
  wire [3:0] _output_instruction_T_6 = input_function7bits[0] ? 4'hc : 4'hb; // @[InstructionChecker.scala 35:12]
  wire [3:0] _output_instruction_T_7 = _output_instruction_T_2 ? _output_instruction_T_4 : _output_instruction_T_6; // @[InstructionChecker.scala 32:26]
  wire [3:0] _output_instruction_T_9 = 7'h3 == input_opcode ? 4'h5 : 4'hf; // @[Mux.scala 81:58]
  wire [3:0] _output_instruction_T_11 = 7'hf == input_opcode ? _output_instruction_T_1 : _output_instruction_T_9; // @[Mux.scala 81:58]
  wire [3:0] _output_instruction_T_13 = 7'h73 == input_opcode ? _output_instruction_T_7 : _output_instruction_T_11; // @[Mux.scala 81:58]
  wire [3:0] _output_instruction_T_15 = 7'h13 == input_opcode ? 4'h7 : _output_instruction_T_13; // @[Mux.scala 81:58]
  wire [3:0] _output_instruction_T_17 = 7'h1b == input_opcode ? 4'h7 : _output_instruction_T_15; // @[Mux.scala 81:58]
  wire [3:0] _output_instruction_T_19 = 7'h67 == input_opcode ? 4'h3 : _output_instruction_T_17; // @[Mux.scala 81:58]
  wire [3:0] _output_instruction_T_21 = 7'h6f == input_opcode ? 4'h2 : _output_instruction_T_19; // @[Mux.scala 81:58]
  wire [3:0] _output_instruction_T_23 = 7'h37 == input_opcode ? 4'h0 : _output_instruction_T_21; // @[Mux.scala 81:58]
  wire [3:0] _output_instruction_T_25 = 7'h17 == input_opcode ? 4'h1 : _output_instruction_T_23; // @[Mux.scala 81:58]
  wire [3:0] _output_instruction_T_27 = 7'h63 == input_opcode ? 4'h4 : _output_instruction_T_25; // @[Mux.scala 81:58]
  wire [3:0] _output_instruction_T_29 = 7'h23 == input_opcode ? 4'h6 : _output_instruction_T_27; // @[Mux.scala 81:58]
  wire [3:0] _output_instruction_T_31 = 7'h33 == input_opcode ? 4'h8 : _output_instruction_T_29; // @[Mux.scala 81:58]
  wire  _output_branch_T = output_instruction == 4'h4; // @[InstructionChecker.scala 56:24]
  wire [2:0] _output_branch_T_2 = 3'h0 == input_function3bits ? 3'h0 : 3'h6; // @[Mux.scala 81:58]
  wire [2:0] _output_branch_T_4 = 3'h1 == input_function3bits ? 3'h1 : _output_branch_T_2; // @[Mux.scala 81:58]
  wire [2:0] _output_branch_T_6 = 3'h4 == input_function3bits ? 3'h2 : _output_branch_T_4; // @[Mux.scala 81:58]
  wire [2:0] _output_branch_T_8 = 3'h5 == input_function3bits ? 3'h3 : _output_branch_T_6; // @[Mux.scala 81:58]
  wire [2:0] _output_branch_T_10 = 3'h6 == input_function3bits ? 3'h4 : _output_branch_T_8; // @[Mux.scala 81:58]
  wire [2:0] _output_branch_T_12 = 3'h7 == input_function3bits ? 3'h5 : _output_branch_T_10; // @[Mux.scala 81:58]
  wire  _output_operationWidth_T_2 = output_instruction == 4'h5 | output_instruction == 4'h6; // @[InstructionChecker.scala 73:46]
  wire [2:0] _output_operationWidth_T_4 = 3'h0 == input_function3bits ? 3'h0 : 3'h4; // @[Mux.scala 81:58]
  wire [2:0] _output_operationWidth_T_6 = 3'h1 == input_function3bits ? 3'h1 : _output_operationWidth_T_4; // @[Mux.scala 81:58]
  wire [2:0] _output_operationWidth_T_8 = 3'h2 == input_function3bits ? 3'h2 : _output_operationWidth_T_6; // @[Mux.scala 81:58]
  wire [2:0] _output_operationWidth_T_10 = 3'h3 == input_function3bits ? 3'h3 : _output_operationWidth_T_8; // @[Mux.scala 81:58]
  wire [6:0] _output_operationWidth_T_11 = input_opcode & 7'h5f; // @[InstructionChecker.scala 87:23]
  wire  _output_operationWidth_T_12 = 7'h13 == _output_operationWidth_T_11; // @[InstructionChecker.scala 87:23]
  wire  _output_operationWidth_T_14 = 7'h1b == _output_operationWidth_T_11; // @[InstructionChecker.scala 88:23]
  wire [2:0] _output_operationWidth_T_15 = _output_operationWidth_T_14 ? 3'h2 : 3'h4; // @[Mux.scala 101:16]
  wire [2:0] _output_operationWidth_T_16 = _output_operationWidth_T_12 ? 3'h3 : _output_operationWidth_T_15; // @[Mux.scala 101:16]
  wire  _output_arithmetic_T = output_instruction == 4'h8; // @[InstructionChecker.scala 94:24]
  wire  _output_arithmetic_T_2 = output_instruction == 4'h8 | output_instruction == 4'h7; // @[InstructionChecker.scala 94:52]
  wire  _output_arithmetic_T_5 = _output_arithmetic_T & input_function7bits[5]; // @[InstructionChecker.scala 100:58]
  wire [2:0] _output_arithmetic_T_8 = input_function7bits[5] ? 3'h7 : 3'h6; // @[InstructionChecker.scala 110:19]
  wire [1:0] _output_arithmetic_T_10 = 3'h1 == input_function3bits ? 2'h2 : {{1'd0}, _output_arithmetic_T_5}; // @[Mux.scala 81:58]
  wire [1:0] _output_arithmetic_T_12 = 3'h2 == input_function3bits ? 2'h3 : _output_arithmetic_T_10; // @[Mux.scala 81:58]
  wire [2:0] _output_arithmetic_T_14 = 3'h3 == input_function3bits ? 3'h4 : {{1'd0}, _output_arithmetic_T_12}; // @[Mux.scala 81:58]
  wire [2:0] _output_arithmetic_T_16 = 3'h4 == input_function3bits ? 3'h5 : _output_arithmetic_T_14; // @[Mux.scala 81:58]
  wire [2:0] _output_arithmetic_T_18 = 3'h5 == input_function3bits ? _output_arithmetic_T_8 : _output_arithmetic_T_16; // @[Mux.scala 81:58]
  wire [3:0] _output_arithmetic_T_20 = 3'h6 == input_function3bits ? 4'h8 : {{1'd0}, _output_arithmetic_T_18}; // @[Mux.scala 81:58]
  wire [3:0] _output_arithmetic_T_22 = 3'h7 == input_function3bits ? 4'h9 : _output_arithmetic_T_20; // @[Mux.scala 81:58]
  assign output_instruction = 7'h3b == input_opcode ? 4'h8 : _output_instruction_T_31; // @[Mux.scala 81:58]
  assign output_branch = _output_branch_T ? _output_branch_T_12 : 3'h6; // @[InstructionChecker.scala 55:23]
  assign output_operationWidth = _output_operationWidth_T_2 ? _output_operationWidth_T_10 : _output_operationWidth_T_16; // @[InstructionChecker.scala 72:31]
  assign output_arithmetic = _output_arithmetic_T_2 ? _output_arithmetic_T_22 : 4'ha; // @[InstructionChecker.scala 93:27]
endmodule
module Executor(
  output        io_reservationStation_ready,
  input         io_reservationStation_valid,
  input         io_reservationStation_bits_destinationTag_threadId,
  input  [3:0]  io_reservationStation_bits_destinationTag_id,
  input  [63:0] io_reservationStation_bits_value1,
  input  [63:0] io_reservationStation_bits_value2,
  input  [2:0]  io_reservationStation_bits_function3,
  input  [11:0] io_reservationStation_bits_immediateOrFunction7,
  input  [6:0]  io_reservationStation_bits_opcode,
  input         io_reservationStation_bits_wasCompressed,
  input         io_out_ready,
  output        io_out_valid,
  output        io_out_bits_resultType,
  output [63:0] io_out_bits_value,
  output        io_out_bits_tag_threadId,
  output [3:0]  io_out_bits_tag_id,
  input         io_fetch_ready,
  output        io_fetch_valid,
  output        io_fetch_bits_threadId,
  output [63:0] io_fetch_bits_programCounterOffset
);
  wire [2:0] instructionChecker_input_function3bits; // @[Executor.scala 31:34]
  wire [6:0] instructionChecker_input_function7bits; // @[Executor.scala 31:34]
  wire [6:0] instructionChecker_input_opcode; // @[Executor.scala 31:34]
  wire [3:0] instructionChecker_output_instruction; // @[Executor.scala 31:34]
  wire [2:0] instructionChecker_output_branch; // @[Executor.scala 31:34]
  wire [2:0] instructionChecker_output_operationWidth; // @[Executor.scala 31:34]
  wire [3:0] instructionChecker_output_arithmetic; // @[Executor.scala 31:34]
  wire [11:0] immediateOrFunction7Extended = io_reservationStation_bits_immediateOrFunction7; // @[Executor.scala 40:53]
  wire [12:0] B_branchedOffset = {io_reservationStation_bits_immediateOrFunction7,1'h0}; // @[Executor.scala 43:55]
  wire  _b_T_1 = instructionChecker_output_instruction == 4'h5; // @[Executor.scala 57:110]
  wire  _b_T_2 = instructionChecker_output_instruction == 4'h7 | instructionChecker_output_instruction == 4'h5; // @[Executor.scala 57:69]
  wire [63:0] b = _b_T_2 ? $signed({{52{immediateOrFunction7Extended[11]}},immediateOrFunction7Extended}) : $signed(
    io_reservationStation_bits_value2); // @[Executor.scala 60:7]
  wire  _executionResult64bit_T = instructionChecker_output_instruction == 4'h6; // @[Executor.scala 66:48]
  wire [63:0] _GEN_10 = {{52{immediateOrFunction7Extended[11]}},immediateOrFunction7Extended}; // @[Executor.scala 66:85]
  wire [63:0] _executionResult64bit_T_4 = $signed(io_reservationStation_bits_value1) + $signed(_GEN_10); // @[Executor.scala 66:85]
  wire [63:0] _executionResult64bit_T_5 = $signed(io_reservationStation_bits_value1) + $signed(_GEN_10); // @[Executor.scala 66:124]
  wire  _executionResult64bit_T_7 = instructionChecker_output_arithmetic == 4'h0; // @[Executor.scala 69:49]
  wire  _executionResult64bit_T_8 = _b_T_1 | _executionResult64bit_T_7; // @[Executor.scala 68:70]
  wire [63:0] _executionResult64bit_T_10 = io_reservationStation_bits_value1 + b; // @[Executor.scala 69:70]
  wire  _executionResult64bit_T_11 = instructionChecker_output_arithmetic == 4'h1; // @[Executor.scala 71:47]
  wire [63:0] _executionResult64bit_T_13 = io_reservationStation_bits_value1 - b; // @[Executor.scala 71:70]
  wire  _executionResult64bit_T_14 = instructionChecker_output_arithmetic == 4'h9; // @[Executor.scala 73:47]
  wire [63:0] _executionResult64bit_T_15 = io_reservationStation_bits_value1 & b; // @[Executor.scala 73:62]
  wire  _executionResult64bit_T_16 = instructionChecker_output_arithmetic == 4'h8; // @[Executor.scala 75:47]
  wire [63:0] _executionResult64bit_T_17 = io_reservationStation_bits_value1 | b; // @[Executor.scala 75:61]
  wire  _executionResult64bit_T_18 = instructionChecker_output_arithmetic == 4'h5; // @[Executor.scala 77:47]
  wire [63:0] _executionResult64bit_T_19 = io_reservationStation_bits_value1 ^ b; // @[Executor.scala 77:62]
  wire  _executionResult64bit_T_20 = instructionChecker_output_arithmetic == 4'h2; // @[Executor.scala 79:47]
  wire  _executionResult64bit_T_21 = instructionChecker_output_operationWidth == 3'h2; // @[Executor.scala 80:52]
  wire [62:0] _GEN_2 = {{31'd0}, io_reservationStation_bits_value1[31:0]}; // @[Executor.scala 81:20]
  wire [62:0] _executionResult64bit_T_24 = _GEN_2 << b[4:0]; // @[Executor.scala 81:20]
  wire [126:0] _GEN_4 = {{63'd0}, io_reservationStation_bits_value1}; // @[Executor.scala 82:13]
  wire [126:0] _executionResult64bit_T_26 = _GEN_4 << b[5:0]; // @[Executor.scala 82:13]
  wire [126:0] _executionResult64bit_T_27 = _executionResult64bit_T_21 ? {{64'd0}, _executionResult64bit_T_24} :
    _executionResult64bit_T_26; // @[Executor.scala 79:75]
  wire  _executionResult64bit_T_28 = instructionChecker_output_arithmetic == 4'h6; // @[Executor.scala 85:47]
  wire [31:0] _executionResult64bit_T_32 = io_reservationStation_bits_value1[31:0] >> b[4:0]; // @[Executor.scala 87:20]
  wire [63:0] _executionResult64bit_T_34 = io_reservationStation_bits_value1 >> b[5:0]; // @[Executor.scala 88:13]
  wire [63:0] _executionResult64bit_T_35 = _executionResult64bit_T_21 ? {{32'd0}, _executionResult64bit_T_32} :
    _executionResult64bit_T_34; // @[Executor.scala 85:97]
  wire  _executionResult64bit_T_36 = instructionChecker_output_arithmetic == 4'h7; // @[Executor.scala 91:47]
  wire [31:0] _executionResult64bit_T_39 = io_reservationStation_bits_value1[31:0]; // @[Executor.scala 93:21]
  wire [31:0] _executionResult64bit_T_42 = $signed(_executionResult64bit_T_39) >>> b[4:0]; // @[Executor.scala 93:40]
  wire [63:0] _executionResult64bit_T_46 = $signed(io_reservationStation_bits_value1) >>> b[5:0]; // @[Executor.scala 94:33]
  wire [63:0] _executionResult64bit_T_47 = _executionResult64bit_T_21 ? {{32'd0}, _executionResult64bit_T_42} :
    _executionResult64bit_T_46; // @[Executor.scala 91:100]
  wire  _executionResult64bit_T_48 = instructionChecker_output_arithmetic == 4'h3; // @[Executor.scala 97:47]
  wire [63:0] _executionResult64bit_T_50 = _b_T_2 ? $signed({{52{immediateOrFunction7Extended[11]}},
    immediateOrFunction7Extended}) : $signed(io_reservationStation_bits_value2); // @[Executor.scala 97:102]
  wire  _executionResult64bit_T_51 = $signed(io_reservationStation_bits_value1) < $signed(_executionResult64bit_T_50); // @[Executor.scala 97:98]
  wire  _executionResult64bit_T_52 = instructionChecker_output_arithmetic == 4'h4; // @[Executor.scala 99:47]
  wire  _executionResult64bit_T_53 = io_reservationStation_bits_value1 < b; // @[Executor.scala 99:99]
  wire  _executionResult64bit_T_55 = instructionChecker_output_instruction == 4'h3; // @[Executor.scala 101:110]
  wire  _executionResult64bit_T_56 = instructionChecker_output_instruction == 4'h2 |
    instructionChecker_output_instruction == 4'h3; // @[Executor.scala 101:69]
  wire [2:0] _executionResult64bit_T_57 = io_reservationStation_bits_wasCompressed ? 3'h2 : 3'h4; // @[Executor.scala 103:16]
  wire [63:0] _GEN_11 = {{61'd0}, _executionResult64bit_T_57}; // @[Executor.scala 102:38]
  wire [63:0] _executionResult64bit_T_59 = io_reservationStation_bits_value2 + _GEN_11; // @[Executor.scala 102:38]
  wire  _executionResult64bit_T_60 = instructionChecker_output_instruction == 4'h0; // @[Executor.scala 105:48]
  wire  _executionResult64bit_T_61 = instructionChecker_output_instruction == 4'h1; // @[Executor.scala 107:48]
  wire [63:0] _executionResult64bit_T_67 = $signed(io_reservationStation_bits_value1) + $signed(
    io_reservationStation_bits_value2); // @[Executor.scala 107:114]
  wire  _executionResult64bit_T_68 = instructionChecker_output_branch == 3'h0; // @[Executor.scala 110:43]
  wire  _executionResult64bit_T_69 = io_reservationStation_bits_value1 == b; // @[Executor.scala 110:77]
  wire  _executionResult64bit_T_70 = instructionChecker_output_branch == 3'h1; // @[Executor.scala 112:43]
  wire  _executionResult64bit_T_71 = io_reservationStation_bits_value1 != b; // @[Executor.scala 112:80]
  wire  _executionResult64bit_T_72 = instructionChecker_output_branch == 3'h2; // @[Executor.scala 114:43]
  wire  _executionResult64bit_T_76 = instructionChecker_output_branch == 3'h4; // @[Executor.scala 116:43]
  wire  _executionResult64bit_T_78 = instructionChecker_output_branch == 3'h3; // @[Executor.scala 118:43]
  wire  _executionResult64bit_T_81 = $signed(io_reservationStation_bits_value1) >= $signed(_executionResult64bit_T_50); // @[Executor.scala 118:93]
  wire  _executionResult64bit_T_82 = instructionChecker_output_branch == 3'h5; // @[Executor.scala 120:43]
  wire  _executionResult64bit_T_83 = io_reservationStation_bits_value1 >= b; // @[Executor.scala 120:94]
  wire  _executionResult64bit_T_85 = _executionResult64bit_T_78 ? _executionResult64bit_T_81 :
    _executionResult64bit_T_82 & _executionResult64bit_T_83; // @[Mux.scala 101:16]
  wire  _executionResult64bit_T_86 = _executionResult64bit_T_76 ? _executionResult64bit_T_53 :
    _executionResult64bit_T_85; // @[Mux.scala 101:16]
  wire  _executionResult64bit_T_87 = _executionResult64bit_T_72 ? _executionResult64bit_T_51 :
    _executionResult64bit_T_86; // @[Mux.scala 101:16]
  wire  _executionResult64bit_T_88 = _executionResult64bit_T_70 ? _executionResult64bit_T_71 :
    _executionResult64bit_T_87; // @[Mux.scala 101:16]
  wire  _executionResult64bit_T_89 = _executionResult64bit_T_68 ? _executionResult64bit_T_69 :
    _executionResult64bit_T_88; // @[Mux.scala 101:16]
  wire [63:0] _executionResult64bit_T_90 = _executionResult64bit_T_61 ? _executionResult64bit_T_67 : {{63'd0},
    _executionResult64bit_T_89}; // @[Mux.scala 101:16]
  wire [63:0] _executionResult64bit_T_91 = _executionResult64bit_T_60 ? io_reservationStation_bits_value1 :
    _executionResult64bit_T_90; // @[Mux.scala 101:16]
  wire [63:0] _executionResult64bit_T_92 = _executionResult64bit_T_56 ? _executionResult64bit_T_59 :
    _executionResult64bit_T_91; // @[Mux.scala 101:16]
  wire [63:0] _executionResult64bit_T_93 = _executionResult64bit_T_52 ? {{63'd0}, _executionResult64bit_T_53} :
    _executionResult64bit_T_92; // @[Mux.scala 101:16]
  wire [63:0] _executionResult64bit_T_94 = _executionResult64bit_T_48 ? {{63'd0}, _executionResult64bit_T_51} :
    _executionResult64bit_T_93; // @[Mux.scala 101:16]
  wire [63:0] _executionResult64bit_T_95 = _executionResult64bit_T_36 ? _executionResult64bit_T_47 :
    _executionResult64bit_T_94; // @[Mux.scala 101:16]
  wire [63:0] _executionResult64bit_T_96 = _executionResult64bit_T_28 ? _executionResult64bit_T_35 :
    _executionResult64bit_T_95; // @[Mux.scala 101:16]
  wire [126:0] _executionResult64bit_T_97 = _executionResult64bit_T_20 ? _executionResult64bit_T_27 : {{63'd0},
    _executionResult64bit_T_96}; // @[Mux.scala 101:16]
  wire [126:0] _executionResult64bit_T_98 = _executionResult64bit_T_18 ? {{63'd0}, _executionResult64bit_T_19} :
    _executionResult64bit_T_97; // @[Mux.scala 101:16]
  wire [126:0] _executionResult64bit_T_99 = _executionResult64bit_T_16 ? {{63'd0}, _executionResult64bit_T_17} :
    _executionResult64bit_T_98; // @[Mux.scala 101:16]
  wire [126:0] _executionResult64bit_T_100 = _executionResult64bit_T_14 ? {{63'd0}, _executionResult64bit_T_15} :
    _executionResult64bit_T_99; // @[Mux.scala 101:16]
  wire [126:0] _executionResult64bit_T_101 = _executionResult64bit_T_11 ? {{63'd0}, _executionResult64bit_T_13} :
    _executionResult64bit_T_100; // @[Mux.scala 101:16]
  wire [126:0] _executionResult64bit_T_102 = _executionResult64bit_T_8 ? {{63'd0}, _executionResult64bit_T_10} :
    _executionResult64bit_T_101; // @[Mux.scala 101:16]
  wire [126:0] _executionResult64bit_T_103 = _executionResult64bit_T ? {{63'd0}, _executionResult64bit_T_5} :
    _executionResult64bit_T_102; // @[Mux.scala 101:16]
  wire [3:0] _io_fetch_bits_programCounterOffset_T = io_reservationStation_bits_wasCompressed ? $signed(4'sh2) :
    $signed(4'sh4); // @[Executor.scala 129:12]
  wire  _io_fetch_bits_programCounterOffset_T_3 = _executionResult64bit_T_68 & _executionResult64bit_T_69; // @[Executor.scala 133:72]
  wire  _io_fetch_bits_programCounterOffset_T_6 = _executionResult64bit_T_70 & _executionResult64bit_T_71; // @[Executor.scala 136:75]
  wire  _io_fetch_bits_programCounterOffset_T_11 = _executionResult64bit_T_72 & _executionResult64bit_T_51; // @[Executor.scala 139:75]
  wire  _io_fetch_bits_programCounterOffset_T_14 = _executionResult64bit_T_76 & _executionResult64bit_T_53; // @[Executor.scala 142:83]
  wire  _io_fetch_bits_programCounterOffset_T_19 = _executionResult64bit_T_78 & _executionResult64bit_T_81; // @[Executor.scala 145:81]
  wire [63:0] _io_fetch_bits_programCounterOffset_T_30 = {_executionResult64bit_T_4[63:1],1'h0}; // @[Executor.scala 155:15]
  wire [63:0] _io_fetch_bits_programCounterOffset_T_34 = $signed(_io_fetch_bits_programCounterOffset_T_30) - $signed(
    io_reservationStation_bits_value2); // @[Executor.scala 155:22]
  wire [63:0] _io_fetch_bits_programCounterOffset_T_35 = _executionResult64bit_T_55 ? $signed(
    _io_fetch_bits_programCounterOffset_T_34) : $signed({{60{_io_fetch_bits_programCounterOffset_T[3]}},
    _io_fetch_bits_programCounterOffset_T}); // @[Mux.scala 101:16]
  wire [63:0] _io_fetch_bits_programCounterOffset_T_36 = _executionResult64bit_T_82 & _executionResult64bit_T_83 ?
    $signed({{51{B_branchedOffset[12]}},B_branchedOffset}) : $signed(_io_fetch_bits_programCounterOffset_T_35); // @[Mux.scala 101:16]
  wire [63:0] _io_fetch_bits_programCounterOffset_T_37 = _io_fetch_bits_programCounterOffset_T_19 ? $signed({{51{
    B_branchedOffset[12]}},B_branchedOffset}) : $signed(_io_fetch_bits_programCounterOffset_T_36); // @[Mux.scala 101:16]
  wire [63:0] _io_fetch_bits_programCounterOffset_T_38 = _io_fetch_bits_programCounterOffset_T_14 ? $signed({{51{
    B_branchedOffset[12]}},B_branchedOffset}) : $signed(_io_fetch_bits_programCounterOffset_T_37); // @[Mux.scala 101:16]
  wire [63:0] _io_fetch_bits_programCounterOffset_T_39 = _io_fetch_bits_programCounterOffset_T_11 ? $signed({{51{
    B_branchedOffset[12]}},B_branchedOffset}) : $signed(_io_fetch_bits_programCounterOffset_T_38); // @[Mux.scala 101:16]
  wire [63:0] _io_fetch_bits_programCounterOffset_T_40 = _io_fetch_bits_programCounterOffset_T_6 ? $signed({{51{
    B_branchedOffset[12]}},B_branchedOffset}) : $signed(_io_fetch_bits_programCounterOffset_T_39); // @[Mux.scala 101:16]
  wire [63:0] _io_fetch_bits_programCounterOffset_T_41 = _io_fetch_bits_programCounterOffset_T_3 ? $signed({{51{
    B_branchedOffset[12]}},B_branchedOffset}) : $signed(_io_fetch_bits_programCounterOffset_T_40); // @[Mux.scala 101:16]
  wire  _GEN_0 = io_fetch_valid & io_reservationStation_bits_destinationTag_threadId; // @[Executor.scala 126:26 127:30 47:26]
  wire [63:0] _GEN_1 = io_fetch_valid ? $signed(_io_fetch_bits_programCounterOffset_T_41) : $signed(64'sh0); // @[Executor.scala 126:26 128:42 45:38]
  wire [126:0] _GEN_3 = io_reservationStation_valid ? _executionResult64bit_T_103 : 127'h0; // @[Executor.scala 49:24 51:37 62:26]
  wire  _executionResultSized_T_3 = ~(_b_T_1 | _executionResult64bit_T); // @[Executor.scala 163:5]
  wire  _executionResultSized_T_5 = _executionResultSized_T_3 & _executionResult64bit_T_21; // @[Executor.scala 165:7]
  wire [63:0] executionResult64bit = _GEN_3[63:0]; // @[Executor.scala 38:34]
  wire [31:0] _executionResultSized_T_7 = executionResult64bit[31:0]; // @[Executor.scala 166:33]
  wire [63:0] _executionResultSized_T_8 = _GEN_3[63:0]; // @[Executor.scala 167:26]
  wire [63:0] executionResultSized = _executionResultSized_T_5 ? $signed({{32{_executionResultSized_T_7[31]}},
    _executionResultSized_T_7}) : $signed(_executionResultSized_T_8); // @[Executor.scala 168:5]
  wire  _io_out_bits_resultType_T = instructionChecker_output_instruction != 4'hf; // @[Executor.scala 179:45]
  wire  _io_out_bits_resultType_T_1 = io_reservationStation_valid & _io_out_bits_resultType_T; // @[Executor.scala 178:33]
  wire  _io_out_bits_resultType_T_2 = instructionChecker_output_instruction != 4'h5; // @[Executor.scala 180:45]
  wire  _io_out_bits_resultType_T_3 = _io_out_bits_resultType_T_1 & _io_out_bits_resultType_T_2; // @[Executor.scala 179:70]
  wire  _io_out_bits_resultType_T_4 = instructionChecker_output_instruction != 4'h6; // @[Executor.scala 181:45]
  wire  _io_out_bits_resultType_T_5 = _io_out_bits_resultType_T_3 & _io_out_bits_resultType_T_4; // @[Executor.scala 180:67]
  InstructionChecker instructionChecker ( // @[Executor.scala 31:34]
    .input_function3bits(instructionChecker_input_function3bits),
    .input_function7bits(instructionChecker_input_function7bits),
    .input_opcode(instructionChecker_input_opcode),
    .output_instruction(instructionChecker_output_instruction),
    .output_branch(instructionChecker_output_branch),
    .output_operationWidth(instructionChecker_output_operationWidth),
    .output_arithmetic(instructionChecker_output_arithmetic)
  );
  assign io_reservationStation_ready = io_out_ready & io_fetch_ready; // @[Executor.scala 30:47]
  assign io_out_valid = io_reservationStation_valid; // @[Executor.scala 48:16 51:37 52:18]
  assign io_out_bits_resultType = _io_out_bits_resultType_T_5 ? 1'h0 : 1'h1; // @[Executor.scala 177:32]
  assign io_out_bits_value = io_out_valid ? executionResultSized : 64'h0; // @[Executor.scala 186:22 188:23 191:23]
  assign io_out_bits_tag_threadId = io_reservationStation_bits_destinationTag_threadId; // @[Executor.scala 186:22 187:21]
  assign io_out_bits_tag_id = io_reservationStation_bits_destinationTag_id; // @[Executor.scala 186:22 187:21]
  assign io_fetch_valid = io_reservationStation_valid & (instructionChecker_output_instruction == 4'h4 |
    _executionResult64bit_T_55); // @[Executor.scala 124:20 46:18 51:37]
  assign io_fetch_bits_threadId = io_reservationStation_valid & _GEN_0; // @[Executor.scala 47:26 51:37]
  assign io_fetch_bits_programCounterOffset = io_reservationStation_valid ? $signed(_GEN_1) : $signed(64'sh0); // @[Executor.scala 51:37 45:38]
  assign instructionChecker_input_function3bits = io_reservationStation_bits_function3; // @[Executor.scala 34:42]
  assign instructionChecker_input_function7bits = io_reservationStation_bits_immediateOrFunction7[11:5]; // @[Executor.scala 36:26]
  assign instructionChecker_input_opcode = io_reservationStation_bits_opcode; // @[Executor.scala 33:35]
endmodule
module Queue_5(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [7:0] io_enq_bits_burstLength,
  input        io_enq_bits_isInstruction,
  input        io_enq_bits_tag_threadId,
  input  [3:0] io_enq_bits_tag_id,
  input  [1:0] io_enq_bits_size,
  input  [2:0] io_enq_bits_offset,
  input        io_enq_bits_signed,
  input        io_deq_ready,
  output       io_deq_valid,
  output [7:0] io_deq_bits_burstLength,
  output       io_deq_bits_isInstruction,
  output       io_deq_bits_tag_threadId,
  output [3:0] io_deq_bits_tag_id,
  output [1:0] io_deq_bits_size,
  output [2:0] io_deq_bits_offset,
  output       io_deq_bits_signed
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_18;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] ram_burstLength [0:7]; // @[Decoupled.scala 273:44]
  wire  ram_burstLength_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:44]
  wire [2:0] ram_burstLength_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:44]
  wire [7:0] ram_burstLength_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:44]
  wire [7:0] ram_burstLength_MPORT_data; // @[Decoupled.scala 273:44]
  wire [2:0] ram_burstLength_MPORT_addr; // @[Decoupled.scala 273:44]
  wire  ram_burstLength_MPORT_mask; // @[Decoupled.scala 273:44]
  wire  ram_burstLength_MPORT_en; // @[Decoupled.scala 273:44]
  reg  ram_burstLength_io_deq_bits_MPORT_en_pipe_0;
  reg [2:0] ram_burstLength_io_deq_bits_MPORT_addr_pipe_0;
  reg  ram_isInstruction [0:7]; // @[Decoupled.scala 273:44]
  wire  ram_isInstruction_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:44]
  wire [2:0] ram_isInstruction_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:44]
  wire  ram_isInstruction_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:44]
  wire  ram_isInstruction_MPORT_data; // @[Decoupled.scala 273:44]
  wire [2:0] ram_isInstruction_MPORT_addr; // @[Decoupled.scala 273:44]
  wire  ram_isInstruction_MPORT_mask; // @[Decoupled.scala 273:44]
  wire  ram_isInstruction_MPORT_en; // @[Decoupled.scala 273:44]
  reg  ram_isInstruction_io_deq_bits_MPORT_en_pipe_0;
  reg [2:0] ram_isInstruction_io_deq_bits_MPORT_addr_pipe_0;
  reg  ram_tag_threadId [0:7]; // @[Decoupled.scala 273:44]
  wire  ram_tag_threadId_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:44]
  wire [2:0] ram_tag_threadId_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:44]
  wire  ram_tag_threadId_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:44]
  wire  ram_tag_threadId_MPORT_data; // @[Decoupled.scala 273:44]
  wire [2:0] ram_tag_threadId_MPORT_addr; // @[Decoupled.scala 273:44]
  wire  ram_tag_threadId_MPORT_mask; // @[Decoupled.scala 273:44]
  wire  ram_tag_threadId_MPORT_en; // @[Decoupled.scala 273:44]
  reg  ram_tag_threadId_io_deq_bits_MPORT_en_pipe_0;
  reg [2:0] ram_tag_threadId_io_deq_bits_MPORT_addr_pipe_0;
  reg [3:0] ram_tag_id [0:7]; // @[Decoupled.scala 273:44]
  wire  ram_tag_id_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:44]
  wire [2:0] ram_tag_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:44]
  wire [3:0] ram_tag_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:44]
  wire [3:0] ram_tag_id_MPORT_data; // @[Decoupled.scala 273:44]
  wire [2:0] ram_tag_id_MPORT_addr; // @[Decoupled.scala 273:44]
  wire  ram_tag_id_MPORT_mask; // @[Decoupled.scala 273:44]
  wire  ram_tag_id_MPORT_en; // @[Decoupled.scala 273:44]
  reg  ram_tag_id_io_deq_bits_MPORT_en_pipe_0;
  reg [2:0] ram_tag_id_io_deq_bits_MPORT_addr_pipe_0;
  reg [1:0] ram_size [0:7]; // @[Decoupled.scala 273:44]
  wire  ram_size_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:44]
  wire [2:0] ram_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:44]
  wire [1:0] ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:44]
  wire [1:0] ram_size_MPORT_data; // @[Decoupled.scala 273:44]
  wire [2:0] ram_size_MPORT_addr; // @[Decoupled.scala 273:44]
  wire  ram_size_MPORT_mask; // @[Decoupled.scala 273:44]
  wire  ram_size_MPORT_en; // @[Decoupled.scala 273:44]
  reg  ram_size_io_deq_bits_MPORT_en_pipe_0;
  reg [2:0] ram_size_io_deq_bits_MPORT_addr_pipe_0;
  reg [2:0] ram_offset [0:7]; // @[Decoupled.scala 273:44]
  wire  ram_offset_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:44]
  wire [2:0] ram_offset_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:44]
  wire [2:0] ram_offset_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:44]
  wire [2:0] ram_offset_MPORT_data; // @[Decoupled.scala 273:44]
  wire [2:0] ram_offset_MPORT_addr; // @[Decoupled.scala 273:44]
  wire  ram_offset_MPORT_mask; // @[Decoupled.scala 273:44]
  wire  ram_offset_MPORT_en; // @[Decoupled.scala 273:44]
  reg  ram_offset_io_deq_bits_MPORT_en_pipe_0;
  reg [2:0] ram_offset_io_deq_bits_MPORT_addr_pipe_0;
  reg  ram_signed [0:7]; // @[Decoupled.scala 273:44]
  wire  ram_signed_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:44]
  wire [2:0] ram_signed_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:44]
  wire  ram_signed_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:44]
  wire  ram_signed_MPORT_data; // @[Decoupled.scala 273:44]
  wire [2:0] ram_signed_MPORT_addr; // @[Decoupled.scala 273:44]
  wire  ram_signed_MPORT_mask; // @[Decoupled.scala 273:44]
  wire  ram_signed_MPORT_en; // @[Decoupled.scala 273:44]
  reg  ram_signed_io_deq_bits_MPORT_en_pipe_0;
  reg [2:0] ram_signed_io_deq_bits_MPORT_addr_pipe_0;
  reg [2:0] enq_ptr_value; // @[Counter.scala 61:40]
  reg [2:0] deq_ptr_value; // @[Counter.scala 61:40]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 277:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 278:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 279:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _value_T_1 = enq_ptr_value + 3'h1; // @[Counter.scala 77:24]
  wire [2:0] _value_T_3 = deq_ptr_value + 3'h1; // @[Counter.scala 77:24]
  wire [3:0] _deq_ptr_next_T_1 = 4'h8 - 4'h1; // @[Decoupled.scala 306:57]
  wire [3:0] _GEN_21 = {{1'd0}, deq_ptr_value}; // @[Decoupled.scala 306:42]
  assign ram_burstLength_io_deq_bits_MPORT_en = ram_burstLength_io_deq_bits_MPORT_en_pipe_0;
  assign ram_burstLength_io_deq_bits_MPORT_addr = ram_burstLength_io_deq_bits_MPORT_addr_pipe_0;
  assign ram_burstLength_io_deq_bits_MPORT_data = ram_burstLength[ram_burstLength_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:44]
  assign ram_burstLength_MPORT_data = io_enq_bits_burstLength;
  assign ram_burstLength_MPORT_addr = enq_ptr_value;
  assign ram_burstLength_MPORT_mask = 1'h1;
  assign ram_burstLength_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_isInstruction_io_deq_bits_MPORT_en = ram_isInstruction_io_deq_bits_MPORT_en_pipe_0;
  assign ram_isInstruction_io_deq_bits_MPORT_addr = ram_isInstruction_io_deq_bits_MPORT_addr_pipe_0;
  assign ram_isInstruction_io_deq_bits_MPORT_data = ram_isInstruction[ram_isInstruction_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:44]
  assign ram_isInstruction_MPORT_data = io_enq_bits_isInstruction;
  assign ram_isInstruction_MPORT_addr = enq_ptr_value;
  assign ram_isInstruction_MPORT_mask = 1'h1;
  assign ram_isInstruction_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_tag_threadId_io_deq_bits_MPORT_en = ram_tag_threadId_io_deq_bits_MPORT_en_pipe_0;
  assign ram_tag_threadId_io_deq_bits_MPORT_addr = ram_tag_threadId_io_deq_bits_MPORT_addr_pipe_0;
  assign ram_tag_threadId_io_deq_bits_MPORT_data = ram_tag_threadId[ram_tag_threadId_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:44]
  assign ram_tag_threadId_MPORT_data = io_enq_bits_tag_threadId;
  assign ram_tag_threadId_MPORT_addr = enq_ptr_value;
  assign ram_tag_threadId_MPORT_mask = 1'h1;
  assign ram_tag_threadId_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_tag_id_io_deq_bits_MPORT_en = ram_tag_id_io_deq_bits_MPORT_en_pipe_0;
  assign ram_tag_id_io_deq_bits_MPORT_addr = ram_tag_id_io_deq_bits_MPORT_addr_pipe_0;
  assign ram_tag_id_io_deq_bits_MPORT_data = ram_tag_id[ram_tag_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:44]
  assign ram_tag_id_MPORT_data = io_enq_bits_tag_id;
  assign ram_tag_id_MPORT_addr = enq_ptr_value;
  assign ram_tag_id_MPORT_mask = 1'h1;
  assign ram_tag_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_size_io_deq_bits_MPORT_en = ram_size_io_deq_bits_MPORT_en_pipe_0;
  assign ram_size_io_deq_bits_MPORT_addr = ram_size_io_deq_bits_MPORT_addr_pipe_0;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:44]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = enq_ptr_value;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_offset_io_deq_bits_MPORT_en = ram_offset_io_deq_bits_MPORT_en_pipe_0;
  assign ram_offset_io_deq_bits_MPORT_addr = ram_offset_io_deq_bits_MPORT_addr_pipe_0;
  assign ram_offset_io_deq_bits_MPORT_data = ram_offset[ram_offset_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:44]
  assign ram_offset_MPORT_data = io_enq_bits_offset;
  assign ram_offset_MPORT_addr = enq_ptr_value;
  assign ram_offset_MPORT_mask = 1'h1;
  assign ram_offset_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_signed_io_deq_bits_MPORT_en = ram_signed_io_deq_bits_MPORT_en_pipe_0;
  assign ram_signed_io_deq_bits_MPORT_addr = ram_signed_io_deq_bits_MPORT_addr_pipe_0;
  assign ram_signed_io_deq_bits_MPORT_data = ram_signed[ram_signed_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:44]
  assign ram_signed_MPORT_data = io_enq_bits_signed;
  assign ram_signed_MPORT_addr = enq_ptr_value;
  assign ram_signed_MPORT_mask = 1'h1;
  assign ram_signed_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 303:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 302:19]
  assign io_deq_bits_burstLength = ram_burstLength_io_deq_bits_MPORT_data; // @[Decoupled.scala 308:17]
  assign io_deq_bits_isInstruction = ram_isInstruction_io_deq_bits_MPORT_data; // @[Decoupled.scala 308:17]
  assign io_deq_bits_tag_threadId = ram_tag_threadId_io_deq_bits_MPORT_data; // @[Decoupled.scala 308:17]
  assign io_deq_bits_tag_id = ram_tag_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 308:17]
  assign io_deq_bits_size = ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 308:17]
  assign io_deq_bits_offset = ram_offset_io_deq_bits_MPORT_data; // @[Decoupled.scala 308:17]
  assign io_deq_bits_signed = ram_signed_io_deq_bits_MPORT_data; // @[Decoupled.scala 308:17]
  always @(posedge clock) begin
    if (ram_burstLength_MPORT_en & ram_burstLength_MPORT_mask) begin
      ram_burstLength[ram_burstLength_MPORT_addr] <= ram_burstLength_MPORT_data; // @[Decoupled.scala 273:44]
    end
    ram_burstLength_io_deq_bits_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (do_deq) begin
        if (_GEN_21 == _deq_ptr_next_T_1) begin // @[Decoupled.scala 306:27]
          ram_burstLength_io_deq_bits_MPORT_addr_pipe_0 <= 3'h0;
        end else begin
          ram_burstLength_io_deq_bits_MPORT_addr_pipe_0 <= _value_T_3;
        end
      end else begin
        ram_burstLength_io_deq_bits_MPORT_addr_pipe_0 <= deq_ptr_value;
      end
    end
    if (ram_isInstruction_MPORT_en & ram_isInstruction_MPORT_mask) begin
      ram_isInstruction[ram_isInstruction_MPORT_addr] <= ram_isInstruction_MPORT_data; // @[Decoupled.scala 273:44]
    end
    ram_isInstruction_io_deq_bits_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (do_deq) begin
        if (_GEN_21 == _deq_ptr_next_T_1) begin // @[Decoupled.scala 306:27]
          ram_isInstruction_io_deq_bits_MPORT_addr_pipe_0 <= 3'h0;
        end else begin
          ram_isInstruction_io_deq_bits_MPORT_addr_pipe_0 <= _value_T_3;
        end
      end else begin
        ram_isInstruction_io_deq_bits_MPORT_addr_pipe_0 <= deq_ptr_value;
      end
    end
    if (ram_tag_threadId_MPORT_en & ram_tag_threadId_MPORT_mask) begin
      ram_tag_threadId[ram_tag_threadId_MPORT_addr] <= ram_tag_threadId_MPORT_data; // @[Decoupled.scala 273:44]
    end
    ram_tag_threadId_io_deq_bits_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (do_deq) begin
        if (_GEN_21 == _deq_ptr_next_T_1) begin // @[Decoupled.scala 306:27]
          ram_tag_threadId_io_deq_bits_MPORT_addr_pipe_0 <= 3'h0;
        end else begin
          ram_tag_threadId_io_deq_bits_MPORT_addr_pipe_0 <= _value_T_3;
        end
      end else begin
        ram_tag_threadId_io_deq_bits_MPORT_addr_pipe_0 <= deq_ptr_value;
      end
    end
    if (ram_tag_id_MPORT_en & ram_tag_id_MPORT_mask) begin
      ram_tag_id[ram_tag_id_MPORT_addr] <= ram_tag_id_MPORT_data; // @[Decoupled.scala 273:44]
    end
    ram_tag_id_io_deq_bits_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (do_deq) begin
        if (_GEN_21 == _deq_ptr_next_T_1) begin // @[Decoupled.scala 306:27]
          ram_tag_id_io_deq_bits_MPORT_addr_pipe_0 <= 3'h0;
        end else begin
          ram_tag_id_io_deq_bits_MPORT_addr_pipe_0 <= _value_T_3;
        end
      end else begin
        ram_tag_id_io_deq_bits_MPORT_addr_pipe_0 <= deq_ptr_value;
      end
    end
    if (ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[Decoupled.scala 273:44]
    end
    ram_size_io_deq_bits_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (do_deq) begin
        if (_GEN_21 == _deq_ptr_next_T_1) begin // @[Decoupled.scala 306:27]
          ram_size_io_deq_bits_MPORT_addr_pipe_0 <= 3'h0;
        end else begin
          ram_size_io_deq_bits_MPORT_addr_pipe_0 <= _value_T_3;
        end
      end else begin
        ram_size_io_deq_bits_MPORT_addr_pipe_0 <= deq_ptr_value;
      end
    end
    if (ram_offset_MPORT_en & ram_offset_MPORT_mask) begin
      ram_offset[ram_offset_MPORT_addr] <= ram_offset_MPORT_data; // @[Decoupled.scala 273:44]
    end
    ram_offset_io_deq_bits_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (do_deq) begin
        if (_GEN_21 == _deq_ptr_next_T_1) begin // @[Decoupled.scala 306:27]
          ram_offset_io_deq_bits_MPORT_addr_pipe_0 <= 3'h0;
        end else begin
          ram_offset_io_deq_bits_MPORT_addr_pipe_0 <= _value_T_3;
        end
      end else begin
        ram_offset_io_deq_bits_MPORT_addr_pipe_0 <= deq_ptr_value;
      end
    end
    if (ram_signed_MPORT_en & ram_signed_MPORT_mask) begin
      ram_signed[ram_signed_MPORT_addr] <= ram_signed_MPORT_data; // @[Decoupled.scala 273:44]
    end
    ram_signed_io_deq_bits_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (do_deq) begin
        if (_GEN_21 == _deq_ptr_next_T_1) begin // @[Decoupled.scala 306:27]
          ram_signed_io_deq_bits_MPORT_addr_pipe_0 <= 3'h0;
        end else begin
          ram_signed_io_deq_bits_MPORT_addr_pipe_0 <= _value_T_3;
        end
      end else begin
        ram_signed_io_deq_bits_MPORT_addr_pipe_0 <= deq_ptr_value;
      end
    end
    if (reset) begin // @[Counter.scala 61:40]
      enq_ptr_value <= 3'h0; // @[Counter.scala 61:40]
    end else if (do_enq) begin // @[Decoupled.scala 286:16]
      enq_ptr_value <= _value_T_1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      deq_ptr_value <= 3'h0; // @[Counter.scala 61:40]
    end else if (do_deq) begin // @[Decoupled.scala 290:16]
      deq_ptr_value <= _value_T_3; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      maybe_full <= do_enq; // @[Decoupled.scala 294:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_burstLength[initvar] = _RAND_0[7:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_isInstruction[initvar] = _RAND_3[0:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_tag_threadId[initvar] = _RAND_6[0:0];
  _RAND_9 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_tag_id[initvar] = _RAND_9[3:0];
  _RAND_12 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_size[initvar] = _RAND_12[1:0];
  _RAND_15 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_offset[initvar] = _RAND_15[2:0];
  _RAND_18 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_signed[initvar] = _RAND_18[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_burstLength_io_deq_bits_MPORT_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  ram_burstLength_io_deq_bits_MPORT_addr_pipe_0 = _RAND_2[2:0];
  _RAND_4 = {1{`RANDOM}};
  ram_isInstruction_io_deq_bits_MPORT_en_pipe_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  ram_isInstruction_io_deq_bits_MPORT_addr_pipe_0 = _RAND_5[2:0];
  _RAND_7 = {1{`RANDOM}};
  ram_tag_threadId_io_deq_bits_MPORT_en_pipe_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  ram_tag_threadId_io_deq_bits_MPORT_addr_pipe_0 = _RAND_8[2:0];
  _RAND_10 = {1{`RANDOM}};
  ram_tag_id_io_deq_bits_MPORT_en_pipe_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  ram_tag_id_io_deq_bits_MPORT_addr_pipe_0 = _RAND_11[2:0];
  _RAND_13 = {1{`RANDOM}};
  ram_size_io_deq_bits_MPORT_en_pipe_0 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  ram_size_io_deq_bits_MPORT_addr_pipe_0 = _RAND_14[2:0];
  _RAND_16 = {1{`RANDOM}};
  ram_offset_io_deq_bits_MPORT_en_pipe_0 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  ram_offset_io_deq_bits_MPORT_addr_pipe_0 = _RAND_17[2:0];
  _RAND_19 = {1{`RANDOM}};
  ram_signed_io_deq_bits_MPORT_en_pipe_0 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  ram_signed_io_deq_bits_MPORT_addr_pipe_0 = _RAND_20[2:0];
  _RAND_21 = {1{`RANDOM}};
  enq_ptr_value = _RAND_21[2:0];
  _RAND_22 = {1{`RANDOM}};
  deq_ptr_value = _RAND_22[2:0];
  _RAND_23 = {1{`RANDOM}};
  maybe_full = _RAND_23[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module FIFO_5(
  input        clock,
  input        reset,
  input        input_valid,
  input  [7:0] input_bits_burstLength,
  input        input_bits_isInstruction,
  input        input_bits_tag_threadId,
  input  [3:0] input_bits_tag_id,
  input  [1:0] input_bits_size,
  input  [2:0] input_bits_offset,
  input        input_bits_signed,
  input        output_ready,
  output [7:0] output_bits_burstLength,
  output       output_bits_isInstruction,
  output       output_bits_tag_threadId,
  output [3:0] output_bits_tag_id,
  output [1:0] output_bits_size,
  output [2:0] output_bits_offset,
  output       output_bits_signed,
  output       full,
  output       empty
);
  wire  queue_clock; // @[FIFO.scala 16:29]
  wire  queue_reset; // @[FIFO.scala 16:29]
  wire  queue_io_enq_ready; // @[FIFO.scala 16:29]
  wire  queue_io_enq_valid; // @[FIFO.scala 16:29]
  wire [7:0] queue_io_enq_bits_burstLength; // @[FIFO.scala 16:29]
  wire  queue_io_enq_bits_isInstruction; // @[FIFO.scala 16:29]
  wire  queue_io_enq_bits_tag_threadId; // @[FIFO.scala 16:29]
  wire [3:0] queue_io_enq_bits_tag_id; // @[FIFO.scala 16:29]
  wire [1:0] queue_io_enq_bits_size; // @[FIFO.scala 16:29]
  wire [2:0] queue_io_enq_bits_offset; // @[FIFO.scala 16:29]
  wire  queue_io_enq_bits_signed; // @[FIFO.scala 16:29]
  wire  queue_io_deq_ready; // @[FIFO.scala 16:29]
  wire  queue_io_deq_valid; // @[FIFO.scala 16:29]
  wire [7:0] queue_io_deq_bits_burstLength; // @[FIFO.scala 16:29]
  wire  queue_io_deq_bits_isInstruction; // @[FIFO.scala 16:29]
  wire  queue_io_deq_bits_tag_threadId; // @[FIFO.scala 16:29]
  wire [3:0] queue_io_deq_bits_tag_id; // @[FIFO.scala 16:29]
  wire [1:0] queue_io_deq_bits_size; // @[FIFO.scala 16:29]
  wire [2:0] queue_io_deq_bits_offset; // @[FIFO.scala 16:29]
  wire  queue_io_deq_bits_signed; // @[FIFO.scala 16:29]
  Queue_5 queue ( // @[FIFO.scala 16:29]
    .clock(queue_clock),
    .reset(queue_reset),
    .io_enq_ready(queue_io_enq_ready),
    .io_enq_valid(queue_io_enq_valid),
    .io_enq_bits_burstLength(queue_io_enq_bits_burstLength),
    .io_enq_bits_isInstruction(queue_io_enq_bits_isInstruction),
    .io_enq_bits_tag_threadId(queue_io_enq_bits_tag_threadId),
    .io_enq_bits_tag_id(queue_io_enq_bits_tag_id),
    .io_enq_bits_size(queue_io_enq_bits_size),
    .io_enq_bits_offset(queue_io_enq_bits_offset),
    .io_enq_bits_signed(queue_io_enq_bits_signed),
    .io_deq_ready(queue_io_deq_ready),
    .io_deq_valid(queue_io_deq_valid),
    .io_deq_bits_burstLength(queue_io_deq_bits_burstLength),
    .io_deq_bits_isInstruction(queue_io_deq_bits_isInstruction),
    .io_deq_bits_tag_threadId(queue_io_deq_bits_tag_threadId),
    .io_deq_bits_tag_id(queue_io_deq_bits_tag_id),
    .io_deq_bits_size(queue_io_deq_bits_size),
    .io_deq_bits_offset(queue_io_deq_bits_offset),
    .io_deq_bits_signed(queue_io_deq_bits_signed)
  );
  assign output_bits_burstLength = queue_io_deq_bits_burstLength; // @[FIFO.scala 20:10]
  assign output_bits_isInstruction = queue_io_deq_bits_isInstruction; // @[FIFO.scala 20:10]
  assign output_bits_tag_threadId = queue_io_deq_bits_tag_threadId; // @[FIFO.scala 20:10]
  assign output_bits_tag_id = queue_io_deq_bits_tag_id; // @[FIFO.scala 20:10]
  assign output_bits_size = queue_io_deq_bits_size; // @[FIFO.scala 20:10]
  assign output_bits_offset = queue_io_deq_bits_offset; // @[FIFO.scala 20:10]
  assign output_bits_signed = queue_io_deq_bits_signed; // @[FIFO.scala 20:10]
  assign full = ~queue_io_enq_ready; // @[FIFO.scala 21:11]
  assign empty = ~queue_io_deq_valid; // @[FIFO.scala 22:12]
  assign queue_clock = clock;
  assign queue_reset = reset;
  assign queue_io_enq_valid = input_valid; // @[FIFO.scala 19:16]
  assign queue_io_enq_bits_burstLength = input_bits_burstLength; // @[FIFO.scala 19:16]
  assign queue_io_enq_bits_isInstruction = input_bits_isInstruction; // @[FIFO.scala 19:16]
  assign queue_io_enq_bits_tag_threadId = input_bits_tag_threadId; // @[FIFO.scala 19:16]
  assign queue_io_enq_bits_tag_id = input_bits_tag_id; // @[FIFO.scala 19:16]
  assign queue_io_enq_bits_size = input_bits_size; // @[FIFO.scala 19:16]
  assign queue_io_enq_bits_offset = input_bits_offset; // @[FIFO.scala 19:16]
  assign queue_io_enq_bits_signed = input_bits_signed; // @[FIFO.scala 19:16]
  assign queue_io_deq_ready = output_ready; // @[FIFO.scala 20:10]
endmodule
module B4RRArbiter_3(
  input         clock,
  input         reset,
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [63:0] io_in_0_bits_address,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [63:0] io_in_1_bits_address,
  input         io_out_ready,
  output        io_out_valid,
  output [63:0] io_out_bits_address,
  output        io_out_bits_outputTag_threadId,
  output        io_chosen
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  _ctrl_validMask_grantMask_lastGrant_T = io_out_ready & io_out_valid; // @[Decoupled.scala 51:35]
  reg  lastGrant; // @[Reg.scala 35:20]
  wire  grantMask_1 = 1'h1 > lastGrant; // @[Arbitar.scala 89:49]
  wire  validMask_1 = io_in_1_valid & grantMask_1; // @[Arbitar.scala 91:57]
  wire  ctrl_2 = ~validMask_1; // @[Arbitar.scala 44:78]
  wire  ctrl_3 = ~(validMask_1 | io_in_0_valid); // @[Arbitar.scala 44:78]
  wire  _T_3 = grantMask_1 | ctrl_3; // @[Arbitar.scala 97:50]
  wire  _GEN_17 = io_in_0_valid ? 1'h0 : 1'h1; // @[Arbitar.scala 102:{26,35} 100:41]
  assign io_in_0_ready = ctrl_2 & io_out_ready; // @[Arbitar.scala 78:21]
  assign io_in_1_ready = _T_3 & io_out_ready; // @[Arbitar.scala 78:21]
  assign io_out_valid = io_chosen ? io_in_1_valid : io_in_0_valid; // @[Arbitar.scala 59:{16,16}]
  assign io_out_bits_address = io_chosen ? io_in_1_bits_address : io_in_0_bits_address; // @[Arbitar.scala 60:{15,15}]
  assign io_out_bits_outputTag_threadId = io_chosen; // @[Arbitar.scala 60:{15,15}]
  assign io_chosen = validMask_1 | _GEN_17; // @[Arbitar.scala 104:{24,33}]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 35:20]
      lastGrant <= 1'h0; // @[Reg.scala 35:20]
    end else if (_ctrl_validMask_grantMask_lastGrant_T) begin // @[Reg.scala 36:18]
      lastGrant <= io_chosen; // @[Reg.scala 36:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  lastGrant = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Arbiter_4(
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [63:0] io_in_0_bits_address,
  input         io_in_0_bits_outputTag_threadId,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [63:0] io_in_1_bits_address,
  input  [1:0]  io_in_1_bits_size,
  input         io_in_1_bits_signed,
  input         io_in_1_bits_outputTag_threadId,
  input  [3:0]  io_in_1_bits_outputTag_id,
  input         io_out_ready,
  output        io_out_valid,
  output        io_out_bits_isInstruction,
  output [63:0] io_out_bits_address,
  output [7:0]  io_out_bits_burstLength,
  output [1:0]  io_out_bits_size,
  output        io_out_bits_signed,
  output        io_out_bits_outputTag_threadId,
  output [3:0]  io_out_bits_outputTag_id
);
  wire  grant_1 = ~io_in_0_valid; // @[Arbiter.scala 45:78]
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 146:19]
  assign io_in_1_ready = grant_1 & io_out_ready; // @[Arbiter.scala 146:19]
  assign io_out_valid = ~grant_1 | io_in_1_valid; // @[Arbiter.scala 147:31]
  assign io_out_bits_isInstruction = io_in_0_valid; // @[Arbiter.scala 136:15 138:26 140:19]
  assign io_out_bits_address = io_in_0_valid ? io_in_0_bits_address : io_in_1_bits_address; // @[Arbiter.scala 136:15 138:26 140:19]
  assign io_out_bits_burstLength = io_in_0_valid ? 8'h1 : 8'h0; // @[Arbiter.scala 136:15 138:26 140:19]
  assign io_out_bits_size = io_in_0_valid ? 2'h3 : io_in_1_bits_size; // @[Arbiter.scala 136:15 138:26 140:19]
  assign io_out_bits_signed = io_in_0_valid ? 1'h0 : io_in_1_bits_signed; // @[Arbiter.scala 136:15 138:26 140:19]
  assign io_out_bits_outputTag_threadId = io_in_0_valid ? io_in_0_bits_outputTag_threadId :
    io_in_1_bits_outputTag_threadId; // @[Arbiter.scala 136:15 138:26 140:19]
  assign io_out_bits_outputTag_id = io_in_0_valid ? 4'h0 : io_in_1_bits_outputTag_id; // @[Arbiter.scala 136:15 138:26 140:19]
endmodule
module Queue_6(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input         io_enq_bits_isInstruction,
  input  [63:0] io_enq_bits_address,
  input  [7:0]  io_enq_bits_burstLength,
  input  [1:0]  io_enq_bits_size,
  input         io_enq_bits_signed,
  input         io_enq_bits_outputTag_threadId,
  input  [3:0]  io_enq_bits_outputTag_id,
  input         io_deq_ready,
  output        io_deq_valid,
  output        io_deq_bits_isInstruction,
  output [63:0] io_deq_bits_address,
  output [7:0]  io_deq_bits_burstLength,
  output [1:0]  io_deq_bits_size,
  output        io_deq_bits_signed,
  output        io_deq_bits_outputTag_threadId,
  output [3:0]  io_deq_bits_outputTag_id
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_18;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
`endif // RANDOMIZE_REG_INIT
  reg  ram_isInstruction [0:3]; // @[Decoupled.scala 273:44]
  wire  ram_isInstruction_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:44]
  wire [1:0] ram_isInstruction_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:44]
  wire  ram_isInstruction_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:44]
  wire  ram_isInstruction_MPORT_data; // @[Decoupled.scala 273:44]
  wire [1:0] ram_isInstruction_MPORT_addr; // @[Decoupled.scala 273:44]
  wire  ram_isInstruction_MPORT_mask; // @[Decoupled.scala 273:44]
  wire  ram_isInstruction_MPORT_en; // @[Decoupled.scala 273:44]
  reg  ram_isInstruction_io_deq_bits_MPORT_en_pipe_0;
  reg [1:0] ram_isInstruction_io_deq_bits_MPORT_addr_pipe_0;
  reg [63:0] ram_address [0:3]; // @[Decoupled.scala 273:44]
  wire  ram_address_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:44]
  wire [1:0] ram_address_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:44]
  wire [63:0] ram_address_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:44]
  wire [63:0] ram_address_MPORT_data; // @[Decoupled.scala 273:44]
  wire [1:0] ram_address_MPORT_addr; // @[Decoupled.scala 273:44]
  wire  ram_address_MPORT_mask; // @[Decoupled.scala 273:44]
  wire  ram_address_MPORT_en; // @[Decoupled.scala 273:44]
  reg  ram_address_io_deq_bits_MPORT_en_pipe_0;
  reg [1:0] ram_address_io_deq_bits_MPORT_addr_pipe_0;
  reg [7:0] ram_burstLength [0:3]; // @[Decoupled.scala 273:44]
  wire  ram_burstLength_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:44]
  wire [1:0] ram_burstLength_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:44]
  wire [7:0] ram_burstLength_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:44]
  wire [7:0] ram_burstLength_MPORT_data; // @[Decoupled.scala 273:44]
  wire [1:0] ram_burstLength_MPORT_addr; // @[Decoupled.scala 273:44]
  wire  ram_burstLength_MPORT_mask; // @[Decoupled.scala 273:44]
  wire  ram_burstLength_MPORT_en; // @[Decoupled.scala 273:44]
  reg  ram_burstLength_io_deq_bits_MPORT_en_pipe_0;
  reg [1:0] ram_burstLength_io_deq_bits_MPORT_addr_pipe_0;
  reg [1:0] ram_size [0:3]; // @[Decoupled.scala 273:44]
  wire  ram_size_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:44]
  wire [1:0] ram_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:44]
  wire [1:0] ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:44]
  wire [1:0] ram_size_MPORT_data; // @[Decoupled.scala 273:44]
  wire [1:0] ram_size_MPORT_addr; // @[Decoupled.scala 273:44]
  wire  ram_size_MPORT_mask; // @[Decoupled.scala 273:44]
  wire  ram_size_MPORT_en; // @[Decoupled.scala 273:44]
  reg  ram_size_io_deq_bits_MPORT_en_pipe_0;
  reg [1:0] ram_size_io_deq_bits_MPORT_addr_pipe_0;
  reg  ram_signed [0:3]; // @[Decoupled.scala 273:44]
  wire  ram_signed_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:44]
  wire [1:0] ram_signed_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:44]
  wire  ram_signed_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:44]
  wire  ram_signed_MPORT_data; // @[Decoupled.scala 273:44]
  wire [1:0] ram_signed_MPORT_addr; // @[Decoupled.scala 273:44]
  wire  ram_signed_MPORT_mask; // @[Decoupled.scala 273:44]
  wire  ram_signed_MPORT_en; // @[Decoupled.scala 273:44]
  reg  ram_signed_io_deq_bits_MPORT_en_pipe_0;
  reg [1:0] ram_signed_io_deq_bits_MPORT_addr_pipe_0;
  reg  ram_outputTag_threadId [0:3]; // @[Decoupled.scala 273:44]
  wire  ram_outputTag_threadId_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:44]
  wire [1:0] ram_outputTag_threadId_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:44]
  wire  ram_outputTag_threadId_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:44]
  wire  ram_outputTag_threadId_MPORT_data; // @[Decoupled.scala 273:44]
  wire [1:0] ram_outputTag_threadId_MPORT_addr; // @[Decoupled.scala 273:44]
  wire  ram_outputTag_threadId_MPORT_mask; // @[Decoupled.scala 273:44]
  wire  ram_outputTag_threadId_MPORT_en; // @[Decoupled.scala 273:44]
  reg  ram_outputTag_threadId_io_deq_bits_MPORT_en_pipe_0;
  reg [1:0] ram_outputTag_threadId_io_deq_bits_MPORT_addr_pipe_0;
  reg [3:0] ram_outputTag_id [0:3]; // @[Decoupled.scala 273:44]
  wire  ram_outputTag_id_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:44]
  wire [1:0] ram_outputTag_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:44]
  wire [3:0] ram_outputTag_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:44]
  wire [3:0] ram_outputTag_id_MPORT_data; // @[Decoupled.scala 273:44]
  wire [1:0] ram_outputTag_id_MPORT_addr; // @[Decoupled.scala 273:44]
  wire  ram_outputTag_id_MPORT_mask; // @[Decoupled.scala 273:44]
  wire  ram_outputTag_id_MPORT_en; // @[Decoupled.scala 273:44]
  reg  ram_outputTag_id_io_deq_bits_MPORT_en_pipe_0;
  reg [1:0] ram_outputTag_id_io_deq_bits_MPORT_addr_pipe_0;
  reg [1:0] enq_ptr_value; // @[Counter.scala 61:40]
  reg [1:0] deq_ptr_value; // @[Counter.scala 61:40]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 277:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 278:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 279:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  wire [1:0] _value_T_1 = enq_ptr_value + 2'h1; // @[Counter.scala 77:24]
  wire [1:0] _value_T_3 = deq_ptr_value + 2'h1; // @[Counter.scala 77:24]
  wire [2:0] _deq_ptr_next_T_1 = 3'h4 - 3'h1; // @[Decoupled.scala 306:57]
  wire [2:0] _GEN_21 = {{1'd0}, deq_ptr_value}; // @[Decoupled.scala 306:42]
  assign ram_isInstruction_io_deq_bits_MPORT_en = ram_isInstruction_io_deq_bits_MPORT_en_pipe_0;
  assign ram_isInstruction_io_deq_bits_MPORT_addr = ram_isInstruction_io_deq_bits_MPORT_addr_pipe_0;
  assign ram_isInstruction_io_deq_bits_MPORT_data = ram_isInstruction[ram_isInstruction_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:44]
  assign ram_isInstruction_MPORT_data = io_enq_bits_isInstruction;
  assign ram_isInstruction_MPORT_addr = enq_ptr_value;
  assign ram_isInstruction_MPORT_mask = 1'h1;
  assign ram_isInstruction_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_address_io_deq_bits_MPORT_en = ram_address_io_deq_bits_MPORT_en_pipe_0;
  assign ram_address_io_deq_bits_MPORT_addr = ram_address_io_deq_bits_MPORT_addr_pipe_0;
  assign ram_address_io_deq_bits_MPORT_data = ram_address[ram_address_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:44]
  assign ram_address_MPORT_data = io_enq_bits_address;
  assign ram_address_MPORT_addr = enq_ptr_value;
  assign ram_address_MPORT_mask = 1'h1;
  assign ram_address_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_burstLength_io_deq_bits_MPORT_en = ram_burstLength_io_deq_bits_MPORT_en_pipe_0;
  assign ram_burstLength_io_deq_bits_MPORT_addr = ram_burstLength_io_deq_bits_MPORT_addr_pipe_0;
  assign ram_burstLength_io_deq_bits_MPORT_data = ram_burstLength[ram_burstLength_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:44]
  assign ram_burstLength_MPORT_data = io_enq_bits_burstLength;
  assign ram_burstLength_MPORT_addr = enq_ptr_value;
  assign ram_burstLength_MPORT_mask = 1'h1;
  assign ram_burstLength_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_size_io_deq_bits_MPORT_en = ram_size_io_deq_bits_MPORT_en_pipe_0;
  assign ram_size_io_deq_bits_MPORT_addr = ram_size_io_deq_bits_MPORT_addr_pipe_0;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:44]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = enq_ptr_value;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_signed_io_deq_bits_MPORT_en = ram_signed_io_deq_bits_MPORT_en_pipe_0;
  assign ram_signed_io_deq_bits_MPORT_addr = ram_signed_io_deq_bits_MPORT_addr_pipe_0;
  assign ram_signed_io_deq_bits_MPORT_data = ram_signed[ram_signed_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:44]
  assign ram_signed_MPORT_data = io_enq_bits_signed;
  assign ram_signed_MPORT_addr = enq_ptr_value;
  assign ram_signed_MPORT_mask = 1'h1;
  assign ram_signed_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_outputTag_threadId_io_deq_bits_MPORT_en = ram_outputTag_threadId_io_deq_bits_MPORT_en_pipe_0;
  assign ram_outputTag_threadId_io_deq_bits_MPORT_addr = ram_outputTag_threadId_io_deq_bits_MPORT_addr_pipe_0;
  assign ram_outputTag_threadId_io_deq_bits_MPORT_data =
    ram_outputTag_threadId[ram_outputTag_threadId_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:44]
  assign ram_outputTag_threadId_MPORT_data = io_enq_bits_outputTag_threadId;
  assign ram_outputTag_threadId_MPORT_addr = enq_ptr_value;
  assign ram_outputTag_threadId_MPORT_mask = 1'h1;
  assign ram_outputTag_threadId_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_outputTag_id_io_deq_bits_MPORT_en = ram_outputTag_id_io_deq_bits_MPORT_en_pipe_0;
  assign ram_outputTag_id_io_deq_bits_MPORT_addr = ram_outputTag_id_io_deq_bits_MPORT_addr_pipe_0;
  assign ram_outputTag_id_io_deq_bits_MPORT_data = ram_outputTag_id[ram_outputTag_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:44]
  assign ram_outputTag_id_MPORT_data = io_enq_bits_outputTag_id;
  assign ram_outputTag_id_MPORT_addr = enq_ptr_value;
  assign ram_outputTag_id_MPORT_mask = 1'h1;
  assign ram_outputTag_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 303:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 302:19]
  assign io_deq_bits_isInstruction = ram_isInstruction_io_deq_bits_MPORT_data; // @[Decoupled.scala 308:17]
  assign io_deq_bits_address = ram_address_io_deq_bits_MPORT_data; // @[Decoupled.scala 308:17]
  assign io_deq_bits_burstLength = ram_burstLength_io_deq_bits_MPORT_data; // @[Decoupled.scala 308:17]
  assign io_deq_bits_size = ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 308:17]
  assign io_deq_bits_signed = ram_signed_io_deq_bits_MPORT_data; // @[Decoupled.scala 308:17]
  assign io_deq_bits_outputTag_threadId = ram_outputTag_threadId_io_deq_bits_MPORT_data; // @[Decoupled.scala 308:17]
  assign io_deq_bits_outputTag_id = ram_outputTag_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 308:17]
  always @(posedge clock) begin
    if (ram_isInstruction_MPORT_en & ram_isInstruction_MPORT_mask) begin
      ram_isInstruction[ram_isInstruction_MPORT_addr] <= ram_isInstruction_MPORT_data; // @[Decoupled.scala 273:44]
    end
    ram_isInstruction_io_deq_bits_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (do_deq) begin
        if (_GEN_21 == _deq_ptr_next_T_1) begin // @[Decoupled.scala 306:27]
          ram_isInstruction_io_deq_bits_MPORT_addr_pipe_0 <= 2'h0;
        end else begin
          ram_isInstruction_io_deq_bits_MPORT_addr_pipe_0 <= _value_T_3;
        end
      end else begin
        ram_isInstruction_io_deq_bits_MPORT_addr_pipe_0 <= deq_ptr_value;
      end
    end
    if (ram_address_MPORT_en & ram_address_MPORT_mask) begin
      ram_address[ram_address_MPORT_addr] <= ram_address_MPORT_data; // @[Decoupled.scala 273:44]
    end
    ram_address_io_deq_bits_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (do_deq) begin
        if (_GEN_21 == _deq_ptr_next_T_1) begin // @[Decoupled.scala 306:27]
          ram_address_io_deq_bits_MPORT_addr_pipe_0 <= 2'h0;
        end else begin
          ram_address_io_deq_bits_MPORT_addr_pipe_0 <= _value_T_3;
        end
      end else begin
        ram_address_io_deq_bits_MPORT_addr_pipe_0 <= deq_ptr_value;
      end
    end
    if (ram_burstLength_MPORT_en & ram_burstLength_MPORT_mask) begin
      ram_burstLength[ram_burstLength_MPORT_addr] <= ram_burstLength_MPORT_data; // @[Decoupled.scala 273:44]
    end
    ram_burstLength_io_deq_bits_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (do_deq) begin
        if (_GEN_21 == _deq_ptr_next_T_1) begin // @[Decoupled.scala 306:27]
          ram_burstLength_io_deq_bits_MPORT_addr_pipe_0 <= 2'h0;
        end else begin
          ram_burstLength_io_deq_bits_MPORT_addr_pipe_0 <= _value_T_3;
        end
      end else begin
        ram_burstLength_io_deq_bits_MPORT_addr_pipe_0 <= deq_ptr_value;
      end
    end
    if (ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[Decoupled.scala 273:44]
    end
    ram_size_io_deq_bits_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (do_deq) begin
        if (_GEN_21 == _deq_ptr_next_T_1) begin // @[Decoupled.scala 306:27]
          ram_size_io_deq_bits_MPORT_addr_pipe_0 <= 2'h0;
        end else begin
          ram_size_io_deq_bits_MPORT_addr_pipe_0 <= _value_T_3;
        end
      end else begin
        ram_size_io_deq_bits_MPORT_addr_pipe_0 <= deq_ptr_value;
      end
    end
    if (ram_signed_MPORT_en & ram_signed_MPORT_mask) begin
      ram_signed[ram_signed_MPORT_addr] <= ram_signed_MPORT_data; // @[Decoupled.scala 273:44]
    end
    ram_signed_io_deq_bits_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (do_deq) begin
        if (_GEN_21 == _deq_ptr_next_T_1) begin // @[Decoupled.scala 306:27]
          ram_signed_io_deq_bits_MPORT_addr_pipe_0 <= 2'h0;
        end else begin
          ram_signed_io_deq_bits_MPORT_addr_pipe_0 <= _value_T_3;
        end
      end else begin
        ram_signed_io_deq_bits_MPORT_addr_pipe_0 <= deq_ptr_value;
      end
    end
    if (ram_outputTag_threadId_MPORT_en & ram_outputTag_threadId_MPORT_mask) begin
      ram_outputTag_threadId[ram_outputTag_threadId_MPORT_addr] <= ram_outputTag_threadId_MPORT_data; // @[Decoupled.scala 273:44]
    end
    ram_outputTag_threadId_io_deq_bits_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (do_deq) begin
        if (_GEN_21 == _deq_ptr_next_T_1) begin // @[Decoupled.scala 306:27]
          ram_outputTag_threadId_io_deq_bits_MPORT_addr_pipe_0 <= 2'h0;
        end else begin
          ram_outputTag_threadId_io_deq_bits_MPORT_addr_pipe_0 <= _value_T_3;
        end
      end else begin
        ram_outputTag_threadId_io_deq_bits_MPORT_addr_pipe_0 <= deq_ptr_value;
      end
    end
    if (ram_outputTag_id_MPORT_en & ram_outputTag_id_MPORT_mask) begin
      ram_outputTag_id[ram_outputTag_id_MPORT_addr] <= ram_outputTag_id_MPORT_data; // @[Decoupled.scala 273:44]
    end
    ram_outputTag_id_io_deq_bits_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (do_deq) begin
        if (_GEN_21 == _deq_ptr_next_T_1) begin // @[Decoupled.scala 306:27]
          ram_outputTag_id_io_deq_bits_MPORT_addr_pipe_0 <= 2'h0;
        end else begin
          ram_outputTag_id_io_deq_bits_MPORT_addr_pipe_0 <= _value_T_3;
        end
      end else begin
        ram_outputTag_id_io_deq_bits_MPORT_addr_pipe_0 <= deq_ptr_value;
      end
    end
    if (reset) begin // @[Counter.scala 61:40]
      enq_ptr_value <= 2'h0; // @[Counter.scala 61:40]
    end else if (do_enq) begin // @[Decoupled.scala 286:16]
      enq_ptr_value <= _value_T_1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      deq_ptr_value <= 2'h0; // @[Counter.scala 61:40]
    end else if (do_deq) begin // @[Decoupled.scala 290:16]
      deq_ptr_value <= _value_T_3; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      maybe_full <= do_enq; // @[Decoupled.scala 294:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_isInstruction[initvar] = _RAND_0[0:0];
  _RAND_3 = {2{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_address[initvar] = _RAND_3[63:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_burstLength[initvar] = _RAND_6[7:0];
  _RAND_9 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_size[initvar] = _RAND_9[1:0];
  _RAND_12 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_signed[initvar] = _RAND_12[0:0];
  _RAND_15 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_outputTag_threadId[initvar] = _RAND_15[0:0];
  _RAND_18 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_outputTag_id[initvar] = _RAND_18[3:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_isInstruction_io_deq_bits_MPORT_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  ram_isInstruction_io_deq_bits_MPORT_addr_pipe_0 = _RAND_2[1:0];
  _RAND_4 = {1{`RANDOM}};
  ram_address_io_deq_bits_MPORT_en_pipe_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  ram_address_io_deq_bits_MPORT_addr_pipe_0 = _RAND_5[1:0];
  _RAND_7 = {1{`RANDOM}};
  ram_burstLength_io_deq_bits_MPORT_en_pipe_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  ram_burstLength_io_deq_bits_MPORT_addr_pipe_0 = _RAND_8[1:0];
  _RAND_10 = {1{`RANDOM}};
  ram_size_io_deq_bits_MPORT_en_pipe_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  ram_size_io_deq_bits_MPORT_addr_pipe_0 = _RAND_11[1:0];
  _RAND_13 = {1{`RANDOM}};
  ram_signed_io_deq_bits_MPORT_en_pipe_0 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  ram_signed_io_deq_bits_MPORT_addr_pipe_0 = _RAND_14[1:0];
  _RAND_16 = {1{`RANDOM}};
  ram_outputTag_threadId_io_deq_bits_MPORT_en_pipe_0 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  ram_outputTag_threadId_io_deq_bits_MPORT_addr_pipe_0 = _RAND_17[1:0];
  _RAND_19 = {1{`RANDOM}};
  ram_outputTag_id_io_deq_bits_MPORT_en_pipe_0 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  ram_outputTag_id_io_deq_bits_MPORT_addr_pipe_0 = _RAND_20[1:0];
  _RAND_21 = {1{`RANDOM}};
  enq_ptr_value = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  deq_ptr_value = _RAND_22[1:0];
  _RAND_23 = {1{`RANDOM}};
  maybe_full = _RAND_23[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module FIFO_6(
  input         clock,
  input         reset,
  output        input_ready,
  input         input_valid,
  input         input_bits_isInstruction,
  input  [63:0] input_bits_address,
  input  [7:0]  input_bits_burstLength,
  input  [1:0]  input_bits_size,
  input         input_bits_signed,
  input         input_bits_outputTag_threadId,
  input  [3:0]  input_bits_outputTag_id,
  input         output_ready,
  output        output_valid,
  output        output_bits_isInstruction,
  output [63:0] output_bits_address,
  output [7:0]  output_bits_burstLength,
  output [1:0]  output_bits_size,
  output        output_bits_signed,
  output        output_bits_outputTag_threadId,
  output [3:0]  output_bits_outputTag_id
);
  wire  queue_clock; // @[FIFO.scala 16:29]
  wire  queue_reset; // @[FIFO.scala 16:29]
  wire  queue_io_enq_ready; // @[FIFO.scala 16:29]
  wire  queue_io_enq_valid; // @[FIFO.scala 16:29]
  wire  queue_io_enq_bits_isInstruction; // @[FIFO.scala 16:29]
  wire [63:0] queue_io_enq_bits_address; // @[FIFO.scala 16:29]
  wire [7:0] queue_io_enq_bits_burstLength; // @[FIFO.scala 16:29]
  wire [1:0] queue_io_enq_bits_size; // @[FIFO.scala 16:29]
  wire  queue_io_enq_bits_signed; // @[FIFO.scala 16:29]
  wire  queue_io_enq_bits_outputTag_threadId; // @[FIFO.scala 16:29]
  wire [3:0] queue_io_enq_bits_outputTag_id; // @[FIFO.scala 16:29]
  wire  queue_io_deq_ready; // @[FIFO.scala 16:29]
  wire  queue_io_deq_valid; // @[FIFO.scala 16:29]
  wire  queue_io_deq_bits_isInstruction; // @[FIFO.scala 16:29]
  wire [63:0] queue_io_deq_bits_address; // @[FIFO.scala 16:29]
  wire [7:0] queue_io_deq_bits_burstLength; // @[FIFO.scala 16:29]
  wire [1:0] queue_io_deq_bits_size; // @[FIFO.scala 16:29]
  wire  queue_io_deq_bits_signed; // @[FIFO.scala 16:29]
  wire  queue_io_deq_bits_outputTag_threadId; // @[FIFO.scala 16:29]
  wire [3:0] queue_io_deq_bits_outputTag_id; // @[FIFO.scala 16:29]
  Queue_6 queue ( // @[FIFO.scala 16:29]
    .clock(queue_clock),
    .reset(queue_reset),
    .io_enq_ready(queue_io_enq_ready),
    .io_enq_valid(queue_io_enq_valid),
    .io_enq_bits_isInstruction(queue_io_enq_bits_isInstruction),
    .io_enq_bits_address(queue_io_enq_bits_address),
    .io_enq_bits_burstLength(queue_io_enq_bits_burstLength),
    .io_enq_bits_size(queue_io_enq_bits_size),
    .io_enq_bits_signed(queue_io_enq_bits_signed),
    .io_enq_bits_outputTag_threadId(queue_io_enq_bits_outputTag_threadId),
    .io_enq_bits_outputTag_id(queue_io_enq_bits_outputTag_id),
    .io_deq_ready(queue_io_deq_ready),
    .io_deq_valid(queue_io_deq_valid),
    .io_deq_bits_isInstruction(queue_io_deq_bits_isInstruction),
    .io_deq_bits_address(queue_io_deq_bits_address),
    .io_deq_bits_burstLength(queue_io_deq_bits_burstLength),
    .io_deq_bits_size(queue_io_deq_bits_size),
    .io_deq_bits_signed(queue_io_deq_bits_signed),
    .io_deq_bits_outputTag_threadId(queue_io_deq_bits_outputTag_threadId),
    .io_deq_bits_outputTag_id(queue_io_deq_bits_outputTag_id)
  );
  assign input_ready = queue_io_enq_ready; // @[FIFO.scala 19:16]
  assign output_valid = queue_io_deq_valid; // @[FIFO.scala 20:10]
  assign output_bits_isInstruction = queue_io_deq_bits_isInstruction; // @[FIFO.scala 20:10]
  assign output_bits_address = queue_io_deq_bits_address; // @[FIFO.scala 20:10]
  assign output_bits_burstLength = queue_io_deq_bits_burstLength; // @[FIFO.scala 20:10]
  assign output_bits_size = queue_io_deq_bits_size; // @[FIFO.scala 20:10]
  assign output_bits_signed = queue_io_deq_bits_signed; // @[FIFO.scala 20:10]
  assign output_bits_outputTag_threadId = queue_io_deq_bits_outputTag_threadId; // @[FIFO.scala 20:10]
  assign output_bits_outputTag_id = queue_io_deq_bits_outputTag_id; // @[FIFO.scala 20:10]
  assign queue_clock = clock;
  assign queue_reset = reset;
  assign queue_io_enq_valid = input_valid; // @[FIFO.scala 19:16]
  assign queue_io_enq_bits_isInstruction = input_bits_isInstruction; // @[FIFO.scala 19:16]
  assign queue_io_enq_bits_address = input_bits_address; // @[FIFO.scala 19:16]
  assign queue_io_enq_bits_burstLength = input_bits_burstLength; // @[FIFO.scala 19:16]
  assign queue_io_enq_bits_size = input_bits_size; // @[FIFO.scala 19:16]
  assign queue_io_enq_bits_signed = input_bits_signed; // @[FIFO.scala 19:16]
  assign queue_io_enq_bits_outputTag_threadId = input_bits_outputTag_threadId; // @[FIFO.scala 19:16]
  assign queue_io_enq_bits_outputTag_id = input_bits_outputTag_id; // @[FIFO.scala 19:16]
  assign queue_io_deq_ready = output_ready; // @[FIFO.scala 20:10]
endmodule
module Queue_7(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [63:0] io_enq_bits_data,
  input  [7:0]  io_enq_bits_strb,
  input         io_deq_ready,
  output        io_deq_valid,
  output [63:0] io_deq_bits_data,
  output [7:0]  io_deq_bits_strb
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] ram_data [0:7]; // @[Decoupled.scala 273:44]
  wire  ram_data_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:44]
  wire [2:0] ram_data_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:44]
  wire [63:0] ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:44]
  wire [63:0] ram_data_MPORT_data; // @[Decoupled.scala 273:44]
  wire [2:0] ram_data_MPORT_addr; // @[Decoupled.scala 273:44]
  wire  ram_data_MPORT_mask; // @[Decoupled.scala 273:44]
  wire  ram_data_MPORT_en; // @[Decoupled.scala 273:44]
  reg  ram_data_io_deq_bits_MPORT_en_pipe_0;
  reg [2:0] ram_data_io_deq_bits_MPORT_addr_pipe_0;
  reg [7:0] ram_strb [0:7]; // @[Decoupled.scala 273:44]
  wire  ram_strb_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:44]
  wire [2:0] ram_strb_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:44]
  wire [7:0] ram_strb_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:44]
  wire [7:0] ram_strb_MPORT_data; // @[Decoupled.scala 273:44]
  wire [2:0] ram_strb_MPORT_addr; // @[Decoupled.scala 273:44]
  wire  ram_strb_MPORT_mask; // @[Decoupled.scala 273:44]
  wire  ram_strb_MPORT_en; // @[Decoupled.scala 273:44]
  reg  ram_strb_io_deq_bits_MPORT_en_pipe_0;
  reg [2:0] ram_strb_io_deq_bits_MPORT_addr_pipe_0;
  reg [2:0] enq_ptr_value; // @[Counter.scala 61:40]
  reg [2:0] deq_ptr_value; // @[Counter.scala 61:40]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 277:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 278:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 279:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _value_T_1 = enq_ptr_value + 3'h1; // @[Counter.scala 77:24]
  wire [2:0] _value_T_3 = deq_ptr_value + 3'h1; // @[Counter.scala 77:24]
  wire [3:0] _deq_ptr_next_T_1 = 4'h8 - 4'h1; // @[Decoupled.scala 306:57]
  wire [3:0] _GEN_16 = {{1'd0}, deq_ptr_value}; // @[Decoupled.scala 306:42]
  assign ram_data_io_deq_bits_MPORT_en = ram_data_io_deq_bits_MPORT_en_pipe_0;
  assign ram_data_io_deq_bits_MPORT_addr = ram_data_io_deq_bits_MPORT_addr_pipe_0;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:44]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = enq_ptr_value;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_strb_io_deq_bits_MPORT_en = ram_strb_io_deq_bits_MPORT_en_pipe_0;
  assign ram_strb_io_deq_bits_MPORT_addr = ram_strb_io_deq_bits_MPORT_addr_pipe_0;
  assign ram_strb_io_deq_bits_MPORT_data = ram_strb[ram_strb_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:44]
  assign ram_strb_MPORT_data = io_enq_bits_strb;
  assign ram_strb_MPORT_addr = enq_ptr_value;
  assign ram_strb_MPORT_mask = 1'h1;
  assign ram_strb_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 303:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 302:19]
  assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 308:17]
  assign io_deq_bits_strb = ram_strb_io_deq_bits_MPORT_data; // @[Decoupled.scala 308:17]
  always @(posedge clock) begin
    if (ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[Decoupled.scala 273:44]
    end
    ram_data_io_deq_bits_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (do_deq) begin
        if (_GEN_16 == _deq_ptr_next_T_1) begin // @[Decoupled.scala 306:27]
          ram_data_io_deq_bits_MPORT_addr_pipe_0 <= 3'h0;
        end else begin
          ram_data_io_deq_bits_MPORT_addr_pipe_0 <= _value_T_3;
        end
      end else begin
        ram_data_io_deq_bits_MPORT_addr_pipe_0 <= deq_ptr_value;
      end
    end
    if (ram_strb_MPORT_en & ram_strb_MPORT_mask) begin
      ram_strb[ram_strb_MPORT_addr] <= ram_strb_MPORT_data; // @[Decoupled.scala 273:44]
    end
    ram_strb_io_deq_bits_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (do_deq) begin
        if (_GEN_16 == _deq_ptr_next_T_1) begin // @[Decoupled.scala 306:27]
          ram_strb_io_deq_bits_MPORT_addr_pipe_0 <= 3'h0;
        end else begin
          ram_strb_io_deq_bits_MPORT_addr_pipe_0 <= _value_T_3;
        end
      end else begin
        ram_strb_io_deq_bits_MPORT_addr_pipe_0 <= deq_ptr_value;
      end
    end
    if (reset) begin // @[Counter.scala 61:40]
      enq_ptr_value <= 3'h0; // @[Counter.scala 61:40]
    end else if (do_enq) begin // @[Decoupled.scala 286:16]
      enq_ptr_value <= _value_T_1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      deq_ptr_value <= 3'h0; // @[Counter.scala 61:40]
    end else if (do_deq) begin // @[Decoupled.scala 290:16]
      deq_ptr_value <= _value_T_3; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      maybe_full <= do_enq; // @[Decoupled.scala 294:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_data[initvar] = _RAND_0[63:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_strb[initvar] = _RAND_3[7:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_data_io_deq_bits_MPORT_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  ram_data_io_deq_bits_MPORT_addr_pipe_0 = _RAND_2[2:0];
  _RAND_4 = {1{`RANDOM}};
  ram_strb_io_deq_bits_MPORT_en_pipe_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  ram_strb_io_deq_bits_MPORT_addr_pipe_0 = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  enq_ptr_value = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  deq_ptr_value = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  maybe_full = _RAND_8[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module FIFO_7(
  input         clock,
  input         reset,
  input         input_valid,
  input  [63:0] input_bits_data,
  input  [7:0]  input_bits_strb,
  input         output_ready,
  output [63:0] output_bits_data,
  output [7:0]  output_bits_strb,
  output        empty
);
  wire  queue_clock; // @[FIFO.scala 16:29]
  wire  queue_reset; // @[FIFO.scala 16:29]
  wire  queue_io_enq_ready; // @[FIFO.scala 16:29]
  wire  queue_io_enq_valid; // @[FIFO.scala 16:29]
  wire [63:0] queue_io_enq_bits_data; // @[FIFO.scala 16:29]
  wire [7:0] queue_io_enq_bits_strb; // @[FIFO.scala 16:29]
  wire  queue_io_deq_ready; // @[FIFO.scala 16:29]
  wire  queue_io_deq_valid; // @[FIFO.scala 16:29]
  wire [63:0] queue_io_deq_bits_data; // @[FIFO.scala 16:29]
  wire [7:0] queue_io_deq_bits_strb; // @[FIFO.scala 16:29]
  Queue_7 queue ( // @[FIFO.scala 16:29]
    .clock(queue_clock),
    .reset(queue_reset),
    .io_enq_ready(queue_io_enq_ready),
    .io_enq_valid(queue_io_enq_valid),
    .io_enq_bits_data(queue_io_enq_bits_data),
    .io_enq_bits_strb(queue_io_enq_bits_strb),
    .io_deq_ready(queue_io_deq_ready),
    .io_deq_valid(queue_io_deq_valid),
    .io_deq_bits_data(queue_io_deq_bits_data),
    .io_deq_bits_strb(queue_io_deq_bits_strb)
  );
  assign output_bits_data = queue_io_deq_bits_data; // @[FIFO.scala 20:10]
  assign output_bits_strb = queue_io_deq_bits_strb; // @[FIFO.scala 20:10]
  assign empty = ~queue_io_deq_valid; // @[FIFO.scala 22:12]
  assign queue_clock = clock;
  assign queue_reset = reset;
  assign queue_io_enq_valid = input_valid; // @[FIFO.scala 19:16]
  assign queue_io_enq_bits_data = input_bits_data; // @[FIFO.scala 19:16]
  assign queue_io_enq_bits_strb = input_bits_strb; // @[FIFO.scala 19:16]
  assign queue_io_deq_ready = output_ready; // @[FIFO.scala 20:10]
endmodule
module Queue_8(
  input   clock,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input   io_deq_ready,
  output  io_deq_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] enq_ptr_value; // @[Counter.scala 61:40]
  reg [2:0] deq_ptr_value; // @[Counter.scala 61:40]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 277:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 278:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 279:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _value_T_1 = enq_ptr_value + 3'h1; // @[Counter.scala 77:24]
  wire [2:0] _value_T_3 = deq_ptr_value + 3'h1; // @[Counter.scala 77:24]
  assign io_enq_ready = ~full; // @[Decoupled.scala 303:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 302:19]
  always @(posedge clock) begin
    if (reset) begin // @[Counter.scala 61:40]
      enq_ptr_value <= 3'h0; // @[Counter.scala 61:40]
    end else if (do_enq) begin // @[Decoupled.scala 286:16]
      enq_ptr_value <= _value_T_1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      deq_ptr_value <= 3'h0; // @[Counter.scala 61:40]
    end else if (do_deq) begin // @[Decoupled.scala 290:16]
      deq_ptr_value <= _value_T_3; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      maybe_full <= do_enq; // @[Decoupled.scala 294:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enq_ptr_value = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  deq_ptr_value = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  maybe_full = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module FIFO_8(
  input   clock,
  input   reset,
  input   input_valid,
  input   output_ready,
  output  empty
);
  wire  queue_clock; // @[FIFO.scala 16:29]
  wire  queue_reset; // @[FIFO.scala 16:29]
  wire  queue_io_enq_ready; // @[FIFO.scala 16:29]
  wire  queue_io_enq_valid; // @[FIFO.scala 16:29]
  wire  queue_io_deq_ready; // @[FIFO.scala 16:29]
  wire  queue_io_deq_valid; // @[FIFO.scala 16:29]
  Queue_8 queue ( // @[FIFO.scala 16:29]
    .clock(queue_clock),
    .reset(queue_reset),
    .io_enq_ready(queue_io_enq_ready),
    .io_enq_valid(queue_io_enq_valid),
    .io_deq_ready(queue_io_deq_ready),
    .io_deq_valid(queue_io_deq_valid)
  );
  assign empty = ~queue_io_deq_valid; // @[FIFO.scala 22:12]
  assign queue_clock = clock;
  assign queue_reset = reset;
  assign queue_io_enq_valid = input_valid; // @[FIFO.scala 19:16]
  assign queue_io_deq_ready = output_ready; // @[FIFO.scala 20:10]
endmodule
module ExternalMemoryInterface(
  input         clock,
  input         reset,
  output        io_dataWriteRequests_ready,
  input         io_dataWriteRequests_valid,
  input  [63:0] io_dataWriteRequests_bits_address,
  input  [63:0] io_dataWriteRequests_bits_data,
  input  [7:0]  io_dataWriteRequests_bits_mask,
  output        io_dataReadRequests_ready,
  input         io_dataReadRequests_valid,
  input  [63:0] io_dataReadRequests_bits_address,
  input  [1:0]  io_dataReadRequests_bits_size,
  input         io_dataReadRequests_bits_signed,
  input         io_dataReadRequests_bits_outputTag_threadId,
  input  [3:0]  io_dataReadRequests_bits_outputTag_id,
  output        io_instructionFetchRequest_0_ready,
  input         io_instructionFetchRequest_0_valid,
  input  [63:0] io_instructionFetchRequest_0_bits_address,
  output        io_instructionFetchRequest_1_ready,
  input         io_instructionFetchRequest_1_valid,
  input  [63:0] io_instructionFetchRequest_1_bits_address,
  input         io_dataReadOut_ready,
  output        io_dataReadOut_valid,
  output [63:0] io_dataReadOut_bits_value,
  output        io_dataReadOut_bits_isError,
  output        io_dataReadOut_bits_tag_threadId,
  output [3:0]  io_dataReadOut_bits_tag_id,
  output        io_instructionOut_0_valid,
  output [63:0] io_instructionOut_0_bits_inner,
  output        io_instructionOut_1_valid,
  output [63:0] io_instructionOut_1_bits_inner,
  input         io_coordinator_writeAddress_ready,
  output        io_coordinator_writeAddress_valid,
  output [63:0] io_coordinator_writeAddress_bits_ADDR,
  output [3:0]  io_coordinator_writeAddress_bits_CACHE,
  input         io_coordinator_write_ready,
  output        io_coordinator_write_valid,
  output [63:0] io_coordinator_write_bits_DATA,
  output [7:0]  io_coordinator_write_bits_STRB,
  output        io_coordinator_write_bits_LAST,
  output        io_coordinator_writeResponse_ready,
  input         io_coordinator_writeResponse_valid,
  input         io_coordinator_readAddress_ready,
  output        io_coordinator_readAddress_valid,
  output [63:0] io_coordinator_readAddress_bits_ADDR,
  output [7:0]  io_coordinator_readAddress_bits_LEN,
  output [3:0]  io_coordinator_readAddress_bits_CACHE,
  output        io_coordinator_read_ready,
  input         io_coordinator_read_valid,
  input  [63:0] io_coordinator_read_bits_DATA,
  input  [1:0]  io_coordinator_read_bits_RESP
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  readQueue_clock; // @[ExternalMemoryInterface.scala 84:25]
  wire  readQueue_reset; // @[ExternalMemoryInterface.scala 84:25]
  wire  readQueue_input_valid; // @[ExternalMemoryInterface.scala 84:25]
  wire [7:0] readQueue_input_bits_burstLength; // @[ExternalMemoryInterface.scala 84:25]
  wire  readQueue_input_bits_isInstruction; // @[ExternalMemoryInterface.scala 84:25]
  wire  readQueue_input_bits_tag_threadId; // @[ExternalMemoryInterface.scala 84:25]
  wire [3:0] readQueue_input_bits_tag_id; // @[ExternalMemoryInterface.scala 84:25]
  wire [1:0] readQueue_input_bits_size; // @[ExternalMemoryInterface.scala 84:25]
  wire [2:0] readQueue_input_bits_offset; // @[ExternalMemoryInterface.scala 84:25]
  wire  readQueue_input_bits_signed; // @[ExternalMemoryInterface.scala 84:25]
  wire  readQueue_output_ready; // @[ExternalMemoryInterface.scala 84:25]
  wire [7:0] readQueue_output_bits_burstLength; // @[ExternalMemoryInterface.scala 84:25]
  wire  readQueue_output_bits_isInstruction; // @[ExternalMemoryInterface.scala 84:25]
  wire  readQueue_output_bits_tag_threadId; // @[ExternalMemoryInterface.scala 84:25]
  wire [3:0] readQueue_output_bits_tag_id; // @[ExternalMemoryInterface.scala 84:25]
  wire [1:0] readQueue_output_bits_size; // @[ExternalMemoryInterface.scala 84:25]
  wire [2:0] readQueue_output_bits_offset; // @[ExternalMemoryInterface.scala 84:25]
  wire  readQueue_output_bits_signed; // @[ExternalMemoryInterface.scala 84:25]
  wire  readQueue_full; // @[ExternalMemoryInterface.scala 84:25]
  wire  readQueue_empty; // @[ExternalMemoryInterface.scala 84:25]
  wire  instructionsArbiter_clock; // @[ExternalMemoryInterface.scala 97:43]
  wire  instructionsArbiter_reset; // @[ExternalMemoryInterface.scala 97:43]
  wire  instructionsArbiter_io_in_0_ready; // @[ExternalMemoryInterface.scala 97:43]
  wire  instructionsArbiter_io_in_0_valid; // @[ExternalMemoryInterface.scala 97:43]
  wire [63:0] instructionsArbiter_io_in_0_bits_address; // @[ExternalMemoryInterface.scala 97:43]
  wire  instructionsArbiter_io_in_1_ready; // @[ExternalMemoryInterface.scala 97:43]
  wire  instructionsArbiter_io_in_1_valid; // @[ExternalMemoryInterface.scala 97:43]
  wire [63:0] instructionsArbiter_io_in_1_bits_address; // @[ExternalMemoryInterface.scala 97:43]
  wire  instructionsArbiter_io_out_ready; // @[ExternalMemoryInterface.scala 97:43]
  wire  instructionsArbiter_io_out_valid; // @[ExternalMemoryInterface.scala 97:43]
  wire [63:0] instructionsArbiter_io_out_bits_address; // @[ExternalMemoryInterface.scala 97:43]
  wire  instructionsArbiter_io_out_bits_outputTag_threadId; // @[ExternalMemoryInterface.scala 97:43]
  wire  instructionsArbiter_io_chosen; // @[ExternalMemoryInterface.scala 97:43]
  wire  instructionOrReadDataArbiter_io_in_0_ready; // @[ExternalMemoryInterface.scala 103:52]
  wire  instructionOrReadDataArbiter_io_in_0_valid; // @[ExternalMemoryInterface.scala 103:52]
  wire [63:0] instructionOrReadDataArbiter_io_in_0_bits_address; // @[ExternalMemoryInterface.scala 103:52]
  wire  instructionOrReadDataArbiter_io_in_0_bits_outputTag_threadId; // @[ExternalMemoryInterface.scala 103:52]
  wire  instructionOrReadDataArbiter_io_in_1_ready; // @[ExternalMemoryInterface.scala 103:52]
  wire  instructionOrReadDataArbiter_io_in_1_valid; // @[ExternalMemoryInterface.scala 103:52]
  wire [63:0] instructionOrReadDataArbiter_io_in_1_bits_address; // @[ExternalMemoryInterface.scala 103:52]
  wire [1:0] instructionOrReadDataArbiter_io_in_1_bits_size; // @[ExternalMemoryInterface.scala 103:52]
  wire  instructionOrReadDataArbiter_io_in_1_bits_signed; // @[ExternalMemoryInterface.scala 103:52]
  wire  instructionOrReadDataArbiter_io_in_1_bits_outputTag_threadId; // @[ExternalMemoryInterface.scala 103:52]
  wire [3:0] instructionOrReadDataArbiter_io_in_1_bits_outputTag_id; // @[ExternalMemoryInterface.scala 103:52]
  wire  instructionOrReadDataArbiter_io_out_ready; // @[ExternalMemoryInterface.scala 103:52]
  wire  instructionOrReadDataArbiter_io_out_valid; // @[ExternalMemoryInterface.scala 103:52]
  wire  instructionOrReadDataArbiter_io_out_bits_isInstruction; // @[ExternalMemoryInterface.scala 103:52]
  wire [63:0] instructionOrReadDataArbiter_io_out_bits_address; // @[ExternalMemoryInterface.scala 103:52]
  wire [7:0] instructionOrReadDataArbiter_io_out_bits_burstLength; // @[ExternalMemoryInterface.scala 103:52]
  wire [1:0] instructionOrReadDataArbiter_io_out_bits_size; // @[ExternalMemoryInterface.scala 103:52]
  wire  instructionOrReadDataArbiter_io_out_bits_signed; // @[ExternalMemoryInterface.scala 103:52]
  wire  instructionOrReadDataArbiter_io_out_bits_outputTag_threadId; // @[ExternalMemoryInterface.scala 103:52]
  wire [3:0] instructionOrReadDataArbiter_io_out_bits_outputTag_id; // @[ExternalMemoryInterface.scala 103:52]
  wire  instructionOrReadDataQueue_clock; // @[ExternalMemoryInterface.scala 108:50]
  wire  instructionOrReadDataQueue_reset; // @[ExternalMemoryInterface.scala 108:50]
  wire  instructionOrReadDataQueue_input_ready; // @[ExternalMemoryInterface.scala 108:50]
  wire  instructionOrReadDataQueue_input_valid; // @[ExternalMemoryInterface.scala 108:50]
  wire  instructionOrReadDataQueue_input_bits_isInstruction; // @[ExternalMemoryInterface.scala 108:50]
  wire [63:0] instructionOrReadDataQueue_input_bits_address; // @[ExternalMemoryInterface.scala 108:50]
  wire [7:0] instructionOrReadDataQueue_input_bits_burstLength; // @[ExternalMemoryInterface.scala 108:50]
  wire [1:0] instructionOrReadDataQueue_input_bits_size; // @[ExternalMemoryInterface.scala 108:50]
  wire  instructionOrReadDataQueue_input_bits_signed; // @[ExternalMemoryInterface.scala 108:50]
  wire  instructionOrReadDataQueue_input_bits_outputTag_threadId; // @[ExternalMemoryInterface.scala 108:50]
  wire [3:0] instructionOrReadDataQueue_input_bits_outputTag_id; // @[ExternalMemoryInterface.scala 108:50]
  wire  instructionOrReadDataQueue_output_ready; // @[ExternalMemoryInterface.scala 108:50]
  wire  instructionOrReadDataQueue_output_valid; // @[ExternalMemoryInterface.scala 108:50]
  wire  instructionOrReadDataQueue_output_bits_isInstruction; // @[ExternalMemoryInterface.scala 108:50]
  wire [63:0] instructionOrReadDataQueue_output_bits_address; // @[ExternalMemoryInterface.scala 108:50]
  wire [7:0] instructionOrReadDataQueue_output_bits_burstLength; // @[ExternalMemoryInterface.scala 108:50]
  wire [1:0] instructionOrReadDataQueue_output_bits_size; // @[ExternalMemoryInterface.scala 108:50]
  wire  instructionOrReadDataQueue_output_bits_signed; // @[ExternalMemoryInterface.scala 108:50]
  wire  instructionOrReadDataQueue_output_bits_outputTag_threadId; // @[ExternalMemoryInterface.scala 108:50]
  wire [3:0] instructionOrReadDataQueue_output_bits_outputTag_id; // @[ExternalMemoryInterface.scala 108:50]
  wire  dataWriteQueue_clock; // @[ExternalMemoryInterface.scala 213:32]
  wire  dataWriteQueue_reset; // @[ExternalMemoryInterface.scala 213:32]
  wire  dataWriteQueue_input_valid; // @[ExternalMemoryInterface.scala 213:32]
  wire [63:0] dataWriteQueue_input_bits_data; // @[ExternalMemoryInterface.scala 213:32]
  wire [7:0] dataWriteQueue_input_bits_strb; // @[ExternalMemoryInterface.scala 213:32]
  wire  dataWriteQueue_output_ready; // @[ExternalMemoryInterface.scala 213:32]
  wire [63:0] dataWriteQueue_output_bits_data; // @[ExternalMemoryInterface.scala 213:32]
  wire [7:0] dataWriteQueue_output_bits_strb; // @[ExternalMemoryInterface.scala 213:32]
  wire  dataWriteQueue_empty; // @[ExternalMemoryInterface.scala 213:32]
  wire  writeResponseQueue_clock; // @[ExternalMemoryInterface.scala 221:36]
  wire  writeResponseQueue_reset; // @[ExternalMemoryInterface.scala 221:36]
  wire  writeResponseQueue_input_valid; // @[ExternalMemoryInterface.scala 221:36]
  wire  writeResponseQueue_output_ready; // @[ExternalMemoryInterface.scala 221:36]
  wire  writeResponseQueue_empty; // @[ExternalMemoryInterface.scala 221:36]
  reg  readQueued; // @[ExternalMemoryInterface.scala 116:27]
  reg [7:0] burstLen; // @[ExternalMemoryInterface.scala 117:25]
  wire [63:0] _io_coordinator_readAddress_bits_ADDR_T_1 = {instructionOrReadDataQueue_output_bits_address[63:3],3'h0}; // @[ExternalMemoryInterface.scala 123:58]
  wire  _GEN_2 = instructionOrReadDataQueue_output_valid; // @[ExternalMemoryInterface.scala 119:33 122:15 48:23]
  wire [63:0] _GEN_3 = instructionOrReadDataQueue_output_valid ? _io_coordinator_readAddress_bits_ADDR_T_1 : 64'h0; // @[ExternalMemoryInterface.scala 119:33 123:19 55:27]
  wire [7:0] _GEN_4 = instructionOrReadDataQueue_output_valid ? instructionOrReadDataQueue_output_bits_burstLength : 8'h0
    ; // @[ExternalMemoryInterface.scala 119:33 124:18 50:26]
  wire [1:0] _GEN_6 = instructionOrReadDataQueue_output_valid ? 2'h2 : 2'h0; // @[ExternalMemoryInterface.scala 119:33 126:20 43:28]
  wire  _GEN_7 = instructionOrReadDataQueue_output_valid & ~readQueued; // @[ExternalMemoryInterface.scala 119:33 128:29 93:25]
  wire  _GEN_16 = instructionOrReadDataQueue_output_valid & io_coordinator_readAddress_ready; // @[ExternalMemoryInterface.scala 114:25 119:33]
  wire  _GEN_17 = readQueue_output_bits_isInstruction | io_dataReadOut_ready; // @[ExternalMemoryInterface.scala 142:49 143:35 145:35]
  wire [7:0] _burstLen_T_1 = burstLen + 8'h1; // @[ExternalMemoryInterface.scala 149:32]
  wire  _T_2 = burstLen == readQueue_output_bits_burstLength; // @[ExternalMemoryInterface.scala 150:25]
  wire [7:0] _GEN_19 = burstLen == readQueue_output_bits_burstLength ? 8'h0 : _burstLen_T_1; // @[ExternalMemoryInterface.scala 149:20 150:64 152:22]
  wire [7:0] _GEN_20 = io_coordinator_read_ready ? _GEN_19 : burstLen; // @[ExternalMemoryInterface.scala 117:25 148:41]
  wire  _GEN_21 = io_coordinator_read_ready & _T_2; // @[ExternalMemoryInterface.scala 148:41 92:26]
  wire  _GEN_22 = ~readQueue_output_bits_tag_threadId; // @[ExternalMemoryInterface.scala 157:{40,40} 79:34]
  wire  _GEN_23 = readQueue_output_bits_tag_threadId; // @[ExternalMemoryInterface.scala 157:{40,40} 79:34]
  wire [63:0] _GEN_24 = ~readQueue_output_bits_tag_threadId ? io_coordinator_read_bits_DATA : 64'h0; // @[ExternalMemoryInterface.scala 159:{45,45} 80:39]
  wire [63:0] _GEN_25 = readQueue_output_bits_tag_threadId ? io_coordinator_read_bits_DATA : 64'h0; // @[ExternalMemoryInterface.scala 159:{45,45} 80:39]
  wire  _io_dataReadOut_bits_value_T = readQueue_output_bits_size == 2'h0; // @[ExternalMemoryInterface.scala 166:43]
  wire  _io_dataReadOut_bits_value_T_1 = readQueue_output_bits_offset == 3'h0; // @[ExternalMemoryInterface.scala 168:49]
  wire  _io_dataReadOut_bits_value_T_3 = readQueue_output_bits_signed & io_coordinator_read_bits_DATA[7]; // @[ExternalMemoryInterface.scala 170:52]
  wire [55:0] _io_dataReadOut_bits_value_T_4 = _io_dataReadOut_bits_value_T_3 ? 56'hffffffffffffff : 56'h0; // @[ExternalMemoryInterface.scala 169:24]
  wire [63:0] _io_dataReadOut_bits_value_T_6 = {_io_dataReadOut_bits_value_T_4,io_coordinator_read_bits_DATA[7:0]}; // @[Cat.scala 33:92]
  wire  _io_dataReadOut_bits_value_T_7 = readQueue_output_bits_offset == 3'h1; // @[ExternalMemoryInterface.scala 168:49]
  wire  _io_dataReadOut_bits_value_T_9 = readQueue_output_bits_signed & io_coordinator_read_bits_DATA[15]; // @[ExternalMemoryInterface.scala 170:52]
  wire [55:0] _io_dataReadOut_bits_value_T_10 = _io_dataReadOut_bits_value_T_9 ? 56'hffffffffffffff : 56'h0; // @[ExternalMemoryInterface.scala 169:24]
  wire [63:0] _io_dataReadOut_bits_value_T_12 = {_io_dataReadOut_bits_value_T_10,io_coordinator_read_bits_DATA[15:8]}; // @[Cat.scala 33:92]
  wire  _io_dataReadOut_bits_value_T_13 = readQueue_output_bits_offset == 3'h2; // @[ExternalMemoryInterface.scala 168:49]
  wire  _io_dataReadOut_bits_value_T_15 = readQueue_output_bits_signed & io_coordinator_read_bits_DATA[23]; // @[ExternalMemoryInterface.scala 170:52]
  wire [55:0] _io_dataReadOut_bits_value_T_16 = _io_dataReadOut_bits_value_T_15 ? 56'hffffffffffffff : 56'h0; // @[ExternalMemoryInterface.scala 169:24]
  wire [63:0] _io_dataReadOut_bits_value_T_18 = {_io_dataReadOut_bits_value_T_16,io_coordinator_read_bits_DATA[23:16]}; // @[Cat.scala 33:92]
  wire  _io_dataReadOut_bits_value_T_19 = readQueue_output_bits_offset == 3'h3; // @[ExternalMemoryInterface.scala 168:49]
  wire  _io_dataReadOut_bits_value_T_21 = readQueue_output_bits_signed & io_coordinator_read_bits_DATA[31]; // @[ExternalMemoryInterface.scala 170:52]
  wire [55:0] _io_dataReadOut_bits_value_T_22 = _io_dataReadOut_bits_value_T_21 ? 56'hffffffffffffff : 56'h0; // @[ExternalMemoryInterface.scala 169:24]
  wire [63:0] _io_dataReadOut_bits_value_T_24 = {_io_dataReadOut_bits_value_T_22,io_coordinator_read_bits_DATA[31:24]}; // @[Cat.scala 33:92]
  wire  _io_dataReadOut_bits_value_T_25 = readQueue_output_bits_offset == 3'h4; // @[ExternalMemoryInterface.scala 168:49]
  wire  _io_dataReadOut_bits_value_T_27 = readQueue_output_bits_signed & io_coordinator_read_bits_DATA[39]; // @[ExternalMemoryInterface.scala 170:52]
  wire [55:0] _io_dataReadOut_bits_value_T_28 = _io_dataReadOut_bits_value_T_27 ? 56'hffffffffffffff : 56'h0; // @[ExternalMemoryInterface.scala 169:24]
  wire [63:0] _io_dataReadOut_bits_value_T_30 = {_io_dataReadOut_bits_value_T_28,io_coordinator_read_bits_DATA[39:32]}; // @[Cat.scala 33:92]
  wire  _io_dataReadOut_bits_value_T_31 = readQueue_output_bits_offset == 3'h5; // @[ExternalMemoryInterface.scala 168:49]
  wire  _io_dataReadOut_bits_value_T_33 = readQueue_output_bits_signed & io_coordinator_read_bits_DATA[47]; // @[ExternalMemoryInterface.scala 170:52]
  wire [55:0] _io_dataReadOut_bits_value_T_34 = _io_dataReadOut_bits_value_T_33 ? 56'hffffffffffffff : 56'h0; // @[ExternalMemoryInterface.scala 169:24]
  wire [63:0] _io_dataReadOut_bits_value_T_36 = {_io_dataReadOut_bits_value_T_34,io_coordinator_read_bits_DATA[47:40]}; // @[Cat.scala 33:92]
  wire  _io_dataReadOut_bits_value_T_37 = readQueue_output_bits_offset == 3'h6; // @[ExternalMemoryInterface.scala 168:49]
  wire  _io_dataReadOut_bits_value_T_39 = readQueue_output_bits_signed & io_coordinator_read_bits_DATA[55]; // @[ExternalMemoryInterface.scala 170:52]
  wire [55:0] _io_dataReadOut_bits_value_T_40 = _io_dataReadOut_bits_value_T_39 ? 56'hffffffffffffff : 56'h0; // @[ExternalMemoryInterface.scala 169:24]
  wire [63:0] _io_dataReadOut_bits_value_T_42 = {_io_dataReadOut_bits_value_T_40,io_coordinator_read_bits_DATA[55:48]}; // @[Cat.scala 33:92]
  wire  _io_dataReadOut_bits_value_T_43 = readQueue_output_bits_offset == 3'h7; // @[ExternalMemoryInterface.scala 168:49]
  wire  _io_dataReadOut_bits_value_T_45 = readQueue_output_bits_signed & io_coordinator_read_bits_DATA[63]; // @[ExternalMemoryInterface.scala 170:52]
  wire [55:0] _io_dataReadOut_bits_value_T_46 = _io_dataReadOut_bits_value_T_45 ? 56'hffffffffffffff : 56'h0; // @[ExternalMemoryInterface.scala 169:24]
  wire [63:0] _io_dataReadOut_bits_value_T_48 = {_io_dataReadOut_bits_value_T_46,io_coordinator_read_bits_DATA[63:56]}; // @[Cat.scala 33:92]
  wire [63:0] _io_dataReadOut_bits_value_T_49 = _io_dataReadOut_bits_value_T_1 ? _io_dataReadOut_bits_value_T_6 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _io_dataReadOut_bits_value_T_50 = _io_dataReadOut_bits_value_T_7 ? _io_dataReadOut_bits_value_T_12 : 64'h0
    ; // @[Mux.scala 27:73]
  wire [63:0] _io_dataReadOut_bits_value_T_51 = _io_dataReadOut_bits_value_T_13 ? _io_dataReadOut_bits_value_T_18 : 64'h0
    ; // @[Mux.scala 27:73]
  wire [63:0] _io_dataReadOut_bits_value_T_52 = _io_dataReadOut_bits_value_T_19 ? _io_dataReadOut_bits_value_T_24 : 64'h0
    ; // @[Mux.scala 27:73]
  wire [63:0] _io_dataReadOut_bits_value_T_53 = _io_dataReadOut_bits_value_T_25 ? _io_dataReadOut_bits_value_T_30 : 64'h0
    ; // @[Mux.scala 27:73]
  wire [63:0] _io_dataReadOut_bits_value_T_54 = _io_dataReadOut_bits_value_T_31 ? _io_dataReadOut_bits_value_T_36 : 64'h0
    ; // @[Mux.scala 27:73]
  wire [63:0] _io_dataReadOut_bits_value_T_55 = _io_dataReadOut_bits_value_T_37 ? _io_dataReadOut_bits_value_T_42 : 64'h0
    ; // @[Mux.scala 27:73]
  wire [63:0] _io_dataReadOut_bits_value_T_56 = _io_dataReadOut_bits_value_T_43 ? _io_dataReadOut_bits_value_T_48 : 64'h0
    ; // @[Mux.scala 27:73]
  wire [63:0] _io_dataReadOut_bits_value_T_57 = _io_dataReadOut_bits_value_T_49 | _io_dataReadOut_bits_value_T_50; // @[Mux.scala 27:73]
  wire [63:0] _io_dataReadOut_bits_value_T_58 = _io_dataReadOut_bits_value_T_57 | _io_dataReadOut_bits_value_T_51; // @[Mux.scala 27:73]
  wire [63:0] _io_dataReadOut_bits_value_T_59 = _io_dataReadOut_bits_value_T_58 | _io_dataReadOut_bits_value_T_52; // @[Mux.scala 27:73]
  wire [63:0] _io_dataReadOut_bits_value_T_60 = _io_dataReadOut_bits_value_T_59 | _io_dataReadOut_bits_value_T_53; // @[Mux.scala 27:73]
  wire [63:0] _io_dataReadOut_bits_value_T_61 = _io_dataReadOut_bits_value_T_60 | _io_dataReadOut_bits_value_T_54; // @[Mux.scala 27:73]
  wire [63:0] _io_dataReadOut_bits_value_T_62 = _io_dataReadOut_bits_value_T_61 | _io_dataReadOut_bits_value_T_55; // @[Mux.scala 27:73]
  wire [63:0] _io_dataReadOut_bits_value_T_63 = _io_dataReadOut_bits_value_T_62 | _io_dataReadOut_bits_value_T_56; // @[Mux.scala 27:73]
  wire  _io_dataReadOut_bits_value_T_64 = readQueue_output_bits_size == 2'h1; // @[ExternalMemoryInterface.scala 178:43]
  wire [47:0] _io_dataReadOut_bits_value_T_68 = _io_dataReadOut_bits_value_T_9 ? 48'hffffffffffff : 48'h0; // @[ExternalMemoryInterface.scala 181:24]
  wire [63:0] _io_dataReadOut_bits_value_T_70 = {_io_dataReadOut_bits_value_T_68,io_coordinator_read_bits_DATA[15:0]}; // @[Cat.scala 33:92]
  wire [47:0] _io_dataReadOut_bits_value_T_74 = _io_dataReadOut_bits_value_T_21 ? 48'hffffffffffff : 48'h0; // @[ExternalMemoryInterface.scala 181:24]
  wire [63:0] _io_dataReadOut_bits_value_T_76 = {_io_dataReadOut_bits_value_T_74,io_coordinator_read_bits_DATA[31:16]}; // @[Cat.scala 33:92]
  wire [47:0] _io_dataReadOut_bits_value_T_80 = _io_dataReadOut_bits_value_T_33 ? 48'hffffffffffff : 48'h0; // @[ExternalMemoryInterface.scala 181:24]
  wire [63:0] _io_dataReadOut_bits_value_T_82 = {_io_dataReadOut_bits_value_T_80,io_coordinator_read_bits_DATA[47:32]}; // @[Cat.scala 33:92]
  wire [47:0] _io_dataReadOut_bits_value_T_86 = _io_dataReadOut_bits_value_T_45 ? 48'hffffffffffff : 48'h0; // @[ExternalMemoryInterface.scala 181:24]
  wire [63:0] _io_dataReadOut_bits_value_T_88 = {_io_dataReadOut_bits_value_T_86,io_coordinator_read_bits_DATA[63:48]}; // @[Cat.scala 33:92]
  wire [63:0] _io_dataReadOut_bits_value_T_89 = _io_dataReadOut_bits_value_T_1 ? _io_dataReadOut_bits_value_T_70 : 64'h0
    ; // @[Mux.scala 27:73]
  wire [63:0] _io_dataReadOut_bits_value_T_90 = _io_dataReadOut_bits_value_T_13 ? _io_dataReadOut_bits_value_T_76 : 64'h0
    ; // @[Mux.scala 27:73]
  wire [63:0] _io_dataReadOut_bits_value_T_91 = _io_dataReadOut_bits_value_T_25 ? _io_dataReadOut_bits_value_T_82 : 64'h0
    ; // @[Mux.scala 27:73]
  wire [63:0] _io_dataReadOut_bits_value_T_92 = _io_dataReadOut_bits_value_T_37 ? _io_dataReadOut_bits_value_T_88 : 64'h0
    ; // @[Mux.scala 27:73]
  wire [63:0] _io_dataReadOut_bits_value_T_93 = _io_dataReadOut_bits_value_T_89 | _io_dataReadOut_bits_value_T_90; // @[Mux.scala 27:73]
  wire [63:0] _io_dataReadOut_bits_value_T_94 = _io_dataReadOut_bits_value_T_93 | _io_dataReadOut_bits_value_T_91; // @[Mux.scala 27:73]
  wire [63:0] _io_dataReadOut_bits_value_T_95 = _io_dataReadOut_bits_value_T_94 | _io_dataReadOut_bits_value_T_92; // @[Mux.scala 27:73]
  wire  _io_dataReadOut_bits_value_T_96 = readQueue_output_bits_size == 2'h2; // @[ExternalMemoryInterface.scala 190:43]
  wire [31:0] _io_dataReadOut_bits_value_T_100 = _io_dataReadOut_bits_value_T_21 ? 32'hffffffff : 32'h0; // @[ExternalMemoryInterface.scala 193:24]
  wire [63:0] _io_dataReadOut_bits_value_T_102 = {_io_dataReadOut_bits_value_T_100,io_coordinator_read_bits_DATA[31:0]}; // @[Cat.scala 33:92]
  wire [31:0] _io_dataReadOut_bits_value_T_106 = _io_dataReadOut_bits_value_T_45 ? 32'hffffffff : 32'h0; // @[ExternalMemoryInterface.scala 193:24]
  wire [63:0] _io_dataReadOut_bits_value_T_108 = {_io_dataReadOut_bits_value_T_106,io_coordinator_read_bits_DATA[63:32]}
    ; // @[Cat.scala 33:92]
  wire [63:0] _io_dataReadOut_bits_value_T_109 = _io_dataReadOut_bits_value_T_1 ? _io_dataReadOut_bits_value_T_102 : 64'h0
    ; // @[Mux.scala 27:73]
  wire [63:0] _io_dataReadOut_bits_value_T_110 = _io_dataReadOut_bits_value_T_25 ? _io_dataReadOut_bits_value_T_108 : 64'h0
    ; // @[Mux.scala 27:73]
  wire [63:0] _io_dataReadOut_bits_value_T_111 = _io_dataReadOut_bits_value_T_109 | _io_dataReadOut_bits_value_T_110; // @[Mux.scala 27:73]
  wire  _io_dataReadOut_bits_value_T_112 = readQueue_output_bits_size == 2'h3; // @[ExternalMemoryInterface.scala 202:43]
  wire [63:0] _io_dataReadOut_bits_value_T_113 = _io_dataReadOut_bits_value_T ? _io_dataReadOut_bits_value_T_63 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _io_dataReadOut_bits_value_T_114 = _io_dataReadOut_bits_value_T_64 ? _io_dataReadOut_bits_value_T_95 : 64'h0
    ; // @[Mux.scala 27:73]
  wire [63:0] _io_dataReadOut_bits_value_T_115 = _io_dataReadOut_bits_value_T_96 ? _io_dataReadOut_bits_value_T_111 : 64'h0
    ; // @[Mux.scala 27:73]
  wire [63:0] _io_dataReadOut_bits_value_T_116 = _io_dataReadOut_bits_value_T_112 ? io_coordinator_read_bits_DATA : 64'h0
    ; // @[Mux.scala 27:73]
  wire [63:0] _io_dataReadOut_bits_value_T_117 = _io_dataReadOut_bits_value_T_113 | _io_dataReadOut_bits_value_T_114; // @[Mux.scala 27:73]
  wire [63:0] _io_dataReadOut_bits_value_T_118 = _io_dataReadOut_bits_value_T_117 | _io_dataReadOut_bits_value_T_115; // @[Mux.scala 27:73]
  wire [63:0] _io_dataReadOut_bits_value_T_119 = _io_dataReadOut_bits_value_T_118 | _io_dataReadOut_bits_value_T_116; // @[Mux.scala 27:73]
  wire  _GEN_26 = readQueue_output_bits_isInstruction & _GEN_22; // @[ExternalMemoryInterface.scala 155:51 79:34]
  wire  _GEN_27 = readQueue_output_bits_isInstruction & _GEN_23; // @[ExternalMemoryInterface.scala 155:51 79:34]
  wire [63:0] _GEN_28 = readQueue_output_bits_isInstruction ? _GEN_24 : 64'h0; // @[ExternalMemoryInterface.scala 155:51 80:39]
  wire [63:0] _GEN_29 = readQueue_output_bits_isInstruction ? _GEN_25 : 64'h0; // @[ExternalMemoryInterface.scala 155:51 80:39]
  wire  _GEN_30 = readQueue_output_bits_isInstruction ? 1'h0 : 1'h1; // @[ExternalMemoryInterface.scala 155:51 76:24 161:32]
  wire  _GEN_31 = readQueue_output_bits_isInstruction ? 1'h0 : readQueue_output_bits_tag_threadId; // @[ExternalMemoryInterface.scala 155:51 72:27 162:35]
  wire [3:0] _GEN_32 = readQueue_output_bits_isInstruction ? 4'h0 : readQueue_output_bits_tag_id; // @[ExternalMemoryInterface.scala 155:51 72:27 162:35]
  wire [63:0] _GEN_33 = readQueue_output_bits_isInstruction ? 64'h0 : _io_dataReadOut_bits_value_T_119; // @[ExternalMemoryInterface.scala 155:51 70:29 164:37]
  wire  _GEN_35 = readQueue_output_bits_isInstruction ? 1'h0 : io_coordinator_read_bits_RESP != 2'h0; // @[ExternalMemoryInterface.scala 155:51 71:31 206:39]
  wire  _GEN_37 = io_coordinator_read_valid & _GEN_21; // @[ExternalMemoryInterface.scala 147:39 92:26]
  wire  _GEN_38 = io_coordinator_read_valid & _GEN_26; // @[ExternalMemoryInterface.scala 147:39 79:34]
  wire  _GEN_39 = io_coordinator_read_valid & _GEN_27; // @[ExternalMemoryInterface.scala 147:39 79:34]
  wire [63:0] _GEN_40 = io_coordinator_read_valid ? _GEN_28 : 64'h0; // @[ExternalMemoryInterface.scala 147:39 80:39]
  wire [63:0] _GEN_41 = io_coordinator_read_valid ? _GEN_29 : 64'h0; // @[ExternalMemoryInterface.scala 147:39 80:39]
  wire  _GEN_42 = io_coordinator_read_valid & _GEN_30; // @[ExternalMemoryInterface.scala 147:39 76:24]
  wire  _GEN_43 = io_coordinator_read_valid & _GEN_31; // @[ExternalMemoryInterface.scala 147:39 72:27]
  wire [3:0] _GEN_44 = io_coordinator_read_valid ? _GEN_32 : 4'h0; // @[ExternalMemoryInterface.scala 147:39 72:27]
  wire [63:0] _GEN_45 = io_coordinator_read_valid ? _GEN_33 : 64'h0; // @[ExternalMemoryInterface.scala 147:39 70:29]
  wire  _GEN_47 = io_coordinator_read_valid & _GEN_35; // @[ExternalMemoryInterface.scala 147:39 71:31]
  wire  _GEN_48 = ~readQueue_empty & _GEN_17; // @[ExternalMemoryInterface.scala 141:28 58:16]
  wire  _GEN_50 = ~readQueue_empty & _GEN_37; // @[ExternalMemoryInterface.scala 141:28 92:26]
  wire  _GEN_51 = ~readQueue_empty & _GEN_38; // @[ExternalMemoryInterface.scala 141:28 79:34]
  wire  _GEN_52 = ~readQueue_empty & _GEN_39; // @[ExternalMemoryInterface.scala 141:28 79:34]
  wire [63:0] _GEN_53 = ~readQueue_empty ? _GEN_40 : 64'h0; // @[ExternalMemoryInterface.scala 141:28 80:39]
  wire [63:0] _GEN_54 = ~readQueue_empty ? _GEN_41 : 64'h0; // @[ExternalMemoryInterface.scala 141:28 80:39]
  wire  _GEN_55 = ~readQueue_empty & _GEN_42; // @[ExternalMemoryInterface.scala 141:28 76:24]
  wire  _GEN_56 = ~readQueue_empty & _GEN_43; // @[ExternalMemoryInterface.scala 141:28 72:27]
  wire [3:0] _GEN_57 = ~readQueue_empty ? _GEN_44 : 4'h0; // @[ExternalMemoryInterface.scala 141:28 72:27]
  wire [63:0] _GEN_58 = ~readQueue_empty ? _GEN_45 : 64'h0; // @[ExternalMemoryInterface.scala 141:28 70:29]
  wire  _GEN_60 = ~readQueue_empty & _GEN_47; // @[ExternalMemoryInterface.scala 141:28 71:31]
  reg  writeQueued; // @[ExternalMemoryInterface.scala 229:30]
  wire  _dataWriteQueue_input_valid_T = ~writeQueued; // @[ExternalMemoryInterface.scala 240:39]
  wire [63:0] _GEN_64 = io_dataWriteRequests_valid ? io_dataWriteRequests_bits_address : 64'h0; // @[ExternalMemoryInterface.scala 230:38 234:19 44:28]
  wire [1:0] _GEN_68 = io_dataWriteRequests_valid ? 2'h2 : 2'h0; // @[ExternalMemoryInterface.scala 230:38 238:20 49:29]
  wire  _GEN_76 = io_dataWriteRequests_valid & io_coordinator_writeAddress_ready; // @[ExternalMemoryInterface.scala 230:38 68:30]
  wire  _T_3 = ~dataWriteQueue_empty; // @[ExternalMemoryInterface.scala 253:10]
  wire [63:0] _GEN_79 = ~dataWriteQueue_empty ? dataWriteQueue_output_bits_data : 64'h0; // @[ExternalMemoryInterface.scala 253:33 255:38 65:21]
  wire [7:0] _GEN_80 = ~dataWriteQueue_empty ? dataWriteQueue_output_bits_strb : 8'h0; // @[ExternalMemoryInterface.scala 253:33 256:38 53:21]
  wire  _T_4 = ~writeResponseQueue_empty; // @[ExternalMemoryInterface.scala 263:10]
  wire [1:0] _GEN_95 = ~readQueue_full ? _GEN_6 : 2'h0; // @[ExternalMemoryInterface.scala 118:25 43:28]
  wire [1:0] _GEN_124 = ~readQueue_full ? _GEN_68 : 2'h0; // @[ExternalMemoryInterface.scala 118:25 49:29]
  FIFO_5 readQueue ( // @[ExternalMemoryInterface.scala 84:25]
    .clock(readQueue_clock),
    .reset(readQueue_reset),
    .input_valid(readQueue_input_valid),
    .input_bits_burstLength(readQueue_input_bits_burstLength),
    .input_bits_isInstruction(readQueue_input_bits_isInstruction),
    .input_bits_tag_threadId(readQueue_input_bits_tag_threadId),
    .input_bits_tag_id(readQueue_input_bits_tag_id),
    .input_bits_size(readQueue_input_bits_size),
    .input_bits_offset(readQueue_input_bits_offset),
    .input_bits_signed(readQueue_input_bits_signed),
    .output_ready(readQueue_output_ready),
    .output_bits_burstLength(readQueue_output_bits_burstLength),
    .output_bits_isInstruction(readQueue_output_bits_isInstruction),
    .output_bits_tag_threadId(readQueue_output_bits_tag_threadId),
    .output_bits_tag_id(readQueue_output_bits_tag_id),
    .output_bits_size(readQueue_output_bits_size),
    .output_bits_offset(readQueue_output_bits_offset),
    .output_bits_signed(readQueue_output_bits_signed),
    .full(readQueue_full),
    .empty(readQueue_empty)
  );
  B4RRArbiter_3 instructionsArbiter ( // @[ExternalMemoryInterface.scala 97:43]
    .clock(instructionsArbiter_clock),
    .reset(instructionsArbiter_reset),
    .io_in_0_ready(instructionsArbiter_io_in_0_ready),
    .io_in_0_valid(instructionsArbiter_io_in_0_valid),
    .io_in_0_bits_address(instructionsArbiter_io_in_0_bits_address),
    .io_in_1_ready(instructionsArbiter_io_in_1_ready),
    .io_in_1_valid(instructionsArbiter_io_in_1_valid),
    .io_in_1_bits_address(instructionsArbiter_io_in_1_bits_address),
    .io_out_ready(instructionsArbiter_io_out_ready),
    .io_out_valid(instructionsArbiter_io_out_valid),
    .io_out_bits_address(instructionsArbiter_io_out_bits_address),
    .io_out_bits_outputTag_threadId(instructionsArbiter_io_out_bits_outputTag_threadId),
    .io_chosen(instructionsArbiter_io_chosen)
  );
  Arbiter_4 instructionOrReadDataArbiter ( // @[ExternalMemoryInterface.scala 103:52]
    .io_in_0_ready(instructionOrReadDataArbiter_io_in_0_ready),
    .io_in_0_valid(instructionOrReadDataArbiter_io_in_0_valid),
    .io_in_0_bits_address(instructionOrReadDataArbiter_io_in_0_bits_address),
    .io_in_0_bits_outputTag_threadId(instructionOrReadDataArbiter_io_in_0_bits_outputTag_threadId),
    .io_in_1_ready(instructionOrReadDataArbiter_io_in_1_ready),
    .io_in_1_valid(instructionOrReadDataArbiter_io_in_1_valid),
    .io_in_1_bits_address(instructionOrReadDataArbiter_io_in_1_bits_address),
    .io_in_1_bits_size(instructionOrReadDataArbiter_io_in_1_bits_size),
    .io_in_1_bits_signed(instructionOrReadDataArbiter_io_in_1_bits_signed),
    .io_in_1_bits_outputTag_threadId(instructionOrReadDataArbiter_io_in_1_bits_outputTag_threadId),
    .io_in_1_bits_outputTag_id(instructionOrReadDataArbiter_io_in_1_bits_outputTag_id),
    .io_out_ready(instructionOrReadDataArbiter_io_out_ready),
    .io_out_valid(instructionOrReadDataArbiter_io_out_valid),
    .io_out_bits_isInstruction(instructionOrReadDataArbiter_io_out_bits_isInstruction),
    .io_out_bits_address(instructionOrReadDataArbiter_io_out_bits_address),
    .io_out_bits_burstLength(instructionOrReadDataArbiter_io_out_bits_burstLength),
    .io_out_bits_size(instructionOrReadDataArbiter_io_out_bits_size),
    .io_out_bits_signed(instructionOrReadDataArbiter_io_out_bits_signed),
    .io_out_bits_outputTag_threadId(instructionOrReadDataArbiter_io_out_bits_outputTag_threadId),
    .io_out_bits_outputTag_id(instructionOrReadDataArbiter_io_out_bits_outputTag_id)
  );
  FIFO_6 instructionOrReadDataQueue ( // @[ExternalMemoryInterface.scala 108:50]
    .clock(instructionOrReadDataQueue_clock),
    .reset(instructionOrReadDataQueue_reset),
    .input_ready(instructionOrReadDataQueue_input_ready),
    .input_valid(instructionOrReadDataQueue_input_valid),
    .input_bits_isInstruction(instructionOrReadDataQueue_input_bits_isInstruction),
    .input_bits_address(instructionOrReadDataQueue_input_bits_address),
    .input_bits_burstLength(instructionOrReadDataQueue_input_bits_burstLength),
    .input_bits_size(instructionOrReadDataQueue_input_bits_size),
    .input_bits_signed(instructionOrReadDataQueue_input_bits_signed),
    .input_bits_outputTag_threadId(instructionOrReadDataQueue_input_bits_outputTag_threadId),
    .input_bits_outputTag_id(instructionOrReadDataQueue_input_bits_outputTag_id),
    .output_ready(instructionOrReadDataQueue_output_ready),
    .output_valid(instructionOrReadDataQueue_output_valid),
    .output_bits_isInstruction(instructionOrReadDataQueue_output_bits_isInstruction),
    .output_bits_address(instructionOrReadDataQueue_output_bits_address),
    .output_bits_burstLength(instructionOrReadDataQueue_output_bits_burstLength),
    .output_bits_size(instructionOrReadDataQueue_output_bits_size),
    .output_bits_signed(instructionOrReadDataQueue_output_bits_signed),
    .output_bits_outputTag_threadId(instructionOrReadDataQueue_output_bits_outputTag_threadId),
    .output_bits_outputTag_id(instructionOrReadDataQueue_output_bits_outputTag_id)
  );
  FIFO_7 dataWriteQueue ( // @[ExternalMemoryInterface.scala 213:32]
    .clock(dataWriteQueue_clock),
    .reset(dataWriteQueue_reset),
    .input_valid(dataWriteQueue_input_valid),
    .input_bits_data(dataWriteQueue_input_bits_data),
    .input_bits_strb(dataWriteQueue_input_bits_strb),
    .output_ready(dataWriteQueue_output_ready),
    .output_bits_data(dataWriteQueue_output_bits_data),
    .output_bits_strb(dataWriteQueue_output_bits_strb),
    .empty(dataWriteQueue_empty)
  );
  FIFO_8 writeResponseQueue ( // @[ExternalMemoryInterface.scala 221:36]
    .clock(writeResponseQueue_clock),
    .reset(writeResponseQueue_reset),
    .input_valid(writeResponseQueue_input_valid),
    .output_ready(writeResponseQueue_output_ready),
    .empty(writeResponseQueue_empty)
  );
  assign io_dataWriteRequests_ready = ~readQueue_full & _GEN_76; // @[ExternalMemoryInterface.scala 118:25 68:30]
  assign io_dataReadRequests_ready = instructionOrReadDataArbiter_io_in_1_ready; // @[ExternalMemoryInterface.scala 107:41]
  assign io_instructionFetchRequest_0_ready = instructionsArbiter_io_in_0_ready; // @[ExternalMemoryInterface.scala 101:36]
  assign io_instructionFetchRequest_1_ready = instructionsArbiter_io_in_1_ready; // @[ExternalMemoryInterface.scala 101:36]
  assign io_dataReadOut_valid = ~readQueue_full & _GEN_55; // @[ExternalMemoryInterface.scala 118:25 76:24]
  assign io_dataReadOut_bits_value = ~readQueue_full ? _GEN_58 : 64'h0; // @[ExternalMemoryInterface.scala 118:25 70:29]
  assign io_dataReadOut_bits_isError = ~readQueue_full & _GEN_60; // @[ExternalMemoryInterface.scala 118:25 71:31]
  assign io_dataReadOut_bits_tag_threadId = ~readQueue_full & _GEN_56; // @[ExternalMemoryInterface.scala 118:25 72:27]
  assign io_dataReadOut_bits_tag_id = ~readQueue_full ? _GEN_57 : 4'h0; // @[ExternalMemoryInterface.scala 118:25 72:27]
  assign io_instructionOut_0_valid = ~readQueue_full & _GEN_51; // @[ExternalMemoryInterface.scala 118:25 79:34]
  assign io_instructionOut_0_bits_inner = ~readQueue_full ? _GEN_53 : 64'h0; // @[ExternalMemoryInterface.scala 118:25 80:39]
  assign io_instructionOut_1_valid = ~readQueue_full & _GEN_52; // @[ExternalMemoryInterface.scala 118:25 79:34]
  assign io_instructionOut_1_bits_inner = ~readQueue_full ? _GEN_54 : 64'h0; // @[ExternalMemoryInterface.scala 118:25 80:39]
  assign io_coordinator_writeAddress_valid = ~readQueue_full & io_dataWriteRequests_valid; // @[ExternalMemoryInterface.scala 118:25 63:24]
  assign io_coordinator_writeAddress_bits_ADDR = ~readQueue_full ? _GEN_64 : 64'h0; // @[ExternalMemoryInterface.scala 118:25 44:28]
  assign io_coordinator_writeAddress_bits_CACHE = {{2'd0}, _GEN_124};
  assign io_coordinator_write_valid = ~readQueue_full & _T_3; // @[ExternalMemoryInterface.scala 118:25 37:17]
  assign io_coordinator_write_bits_DATA = ~readQueue_full ? _GEN_79 : 64'h0; // @[ExternalMemoryInterface.scala 118:25 65:21]
  assign io_coordinator_write_bits_STRB = ~readQueue_full ? _GEN_80 : 8'h0; // @[ExternalMemoryInterface.scala 118:25 53:21]
  assign io_coordinator_write_bits_LAST = ~readQueue_full & _T_3; // @[ExternalMemoryInterface.scala 118:25 37:17]
  assign io_coordinator_writeResponse_ready = ~readQueue_full & _T_4; // @[ExternalMemoryInterface.scala 118:25 36:25]
  assign io_coordinator_readAddress_valid = ~readQueue_full & _GEN_2; // @[ExternalMemoryInterface.scala 118:25 48:23]
  assign io_coordinator_readAddress_bits_ADDR = ~readQueue_full ? _GEN_3 : 64'h0; // @[ExternalMemoryInterface.scala 118:25 55:27]
  assign io_coordinator_readAddress_bits_LEN = ~readQueue_full ? _GEN_4 : 8'h0; // @[ExternalMemoryInterface.scala 118:25 50:26]
  assign io_coordinator_readAddress_bits_CACHE = {{2'd0}, _GEN_95};
  assign io_coordinator_read_ready = ~readQueue_full & _GEN_48; // @[ExternalMemoryInterface.scala 118:25 58:16]
  assign readQueue_clock = clock;
  assign readQueue_reset = reset;
  assign readQueue_input_valid = ~readQueue_full & _GEN_7; // @[ExternalMemoryInterface.scala 118:25 93:25]
  assign readQueue_input_bits_burstLength = instructionOrReadDataQueue_output_bits_burstLength; // @[ExternalMemoryInterface.scala 119:33 129:40]
  assign readQueue_input_bits_isInstruction = instructionOrReadDataQueue_output_bits_isInstruction; // @[ExternalMemoryInterface.scala 119:33 130:42]
  assign readQueue_input_bits_tag_threadId = instructionOrReadDataQueue_output_bits_outputTag_threadId; // @[ExternalMemoryInterface.scala 119:33 131:32]
  assign readQueue_input_bits_tag_id = instructionOrReadDataQueue_output_bits_outputTag_id; // @[ExternalMemoryInterface.scala 119:33 131:32]
  assign readQueue_input_bits_size = instructionOrReadDataQueue_output_bits_size; // @[ExternalMemoryInterface.scala 119:33 133:33]
  assign readQueue_input_bits_offset = instructionOrReadDataQueue_output_bits_address[2:0]; // @[ExternalMemoryInterface.scala 132:66]
  assign readQueue_input_bits_signed = instructionOrReadDataQueue_output_bits_signed; // @[ExternalMemoryInterface.scala 119:33 134:35]
  assign readQueue_output_ready = ~readQueue_full & _GEN_50; // @[ExternalMemoryInterface.scala 118:25 92:26]
  assign instructionsArbiter_clock = clock;
  assign instructionsArbiter_reset = reset;
  assign instructionsArbiter_io_in_0_valid = io_instructionFetchRequest_0_valid; // @[ExternalMemoryInterface.scala 101:36]
  assign instructionsArbiter_io_in_0_bits_address = io_instructionFetchRequest_0_bits_address; // @[ExternalMemoryInterface.scala 101:36]
  assign instructionsArbiter_io_in_1_valid = io_instructionFetchRequest_1_valid; // @[ExternalMemoryInterface.scala 101:36]
  assign instructionsArbiter_io_in_1_bits_address = io_instructionFetchRequest_1_bits_address; // @[ExternalMemoryInterface.scala 101:36]
  assign instructionsArbiter_io_out_ready = instructionOrReadDataArbiter_io_in_0_ready; // @[ExternalMemoryInterface.scala 106:41]
  assign instructionOrReadDataArbiter_io_in_0_valid = instructionsArbiter_io_out_valid; // @[ExternalMemoryInterface.scala 106:41]
  assign instructionOrReadDataArbiter_io_in_0_bits_address = instructionsArbiter_io_out_bits_address; // @[ExternalMemoryInterface.scala 106:41]
  assign instructionOrReadDataArbiter_io_in_0_bits_outputTag_threadId =
    instructionsArbiter_io_out_bits_outputTag_threadId; // @[ExternalMemoryInterface.scala 106:41]
  assign instructionOrReadDataArbiter_io_in_1_valid = io_dataReadRequests_valid; // @[ExternalMemoryInterface.scala 107:41]
  assign instructionOrReadDataArbiter_io_in_1_bits_address = io_dataReadRequests_bits_address; // @[ExternalMemoryInterface.scala 107:41]
  assign instructionOrReadDataArbiter_io_in_1_bits_size = io_dataReadRequests_bits_size; // @[ExternalMemoryInterface.scala 107:41]
  assign instructionOrReadDataArbiter_io_in_1_bits_signed = io_dataReadRequests_bits_signed; // @[ExternalMemoryInterface.scala 107:41]
  assign instructionOrReadDataArbiter_io_in_1_bits_outputTag_threadId = io_dataReadRequests_bits_outputTag_threadId; // @[ExternalMemoryInterface.scala 107:41]
  assign instructionOrReadDataArbiter_io_in_1_bits_outputTag_id = io_dataReadRequests_bits_outputTag_id; // @[ExternalMemoryInterface.scala 107:41]
  assign instructionOrReadDataArbiter_io_out_ready = instructionOrReadDataQueue_input_ready; // @[ExternalMemoryInterface.scala 111:36]
  assign instructionOrReadDataQueue_clock = clock;
  assign instructionOrReadDataQueue_reset = reset;
  assign instructionOrReadDataQueue_input_valid = instructionOrReadDataArbiter_io_out_valid; // @[ExternalMemoryInterface.scala 111:36]
  assign instructionOrReadDataQueue_input_bits_isInstruction = instructionOrReadDataArbiter_io_out_bits_isInstruction; // @[ExternalMemoryInterface.scala 111:36]
  assign instructionOrReadDataQueue_input_bits_address = instructionOrReadDataArbiter_io_out_bits_address; // @[ExternalMemoryInterface.scala 111:36]
  assign instructionOrReadDataQueue_input_bits_burstLength = instructionOrReadDataArbiter_io_out_bits_burstLength; // @[ExternalMemoryInterface.scala 111:36]
  assign instructionOrReadDataQueue_input_bits_size = instructionOrReadDataArbiter_io_out_bits_size; // @[ExternalMemoryInterface.scala 111:36]
  assign instructionOrReadDataQueue_input_bits_signed = instructionOrReadDataArbiter_io_out_bits_signed; // @[ExternalMemoryInterface.scala 111:36]
  assign instructionOrReadDataQueue_input_bits_outputTag_threadId =
    instructionOrReadDataArbiter_io_out_bits_outputTag_threadId; // @[ExternalMemoryInterface.scala 111:36]
  assign instructionOrReadDataQueue_input_bits_outputTag_id = instructionOrReadDataArbiter_io_out_bits_outputTag_id; // @[ExternalMemoryInterface.scala 111:36]
  assign instructionOrReadDataQueue_output_ready = ~readQueue_full & _GEN_16; // @[ExternalMemoryInterface.scala 114:25 118:25]
  assign dataWriteQueue_clock = clock;
  assign dataWriteQueue_reset = reset;
  assign dataWriteQueue_input_valid = io_dataWriteRequests_valid & ~writeQueued; // @[ExternalMemoryInterface.scala 218:32 230:38 240:36]
  assign dataWriteQueue_input_bits_data = io_dataWriteRequests_bits_data; // @[ExternalMemoryInterface.scala 230:38 241:40]
  assign dataWriteQueue_input_bits_strb = io_dataWriteRequests_bits_mask; // @[ExternalMemoryInterface.scala 230:38 242:40]
  assign dataWriteQueue_output_ready = ~dataWriteQueue_empty & io_coordinator_write_ready; // @[ExternalMemoryInterface.scala 217:33 253:33]
  assign writeResponseQueue_clock = clock;
  assign writeResponseQueue_reset = reset;
  assign writeResponseQueue_input_valid = io_dataWriteRequests_valid & _dataWriteQueue_input_valid_T; // @[ExternalMemoryInterface.scala 225:36 230:38 243:40]
  assign writeResponseQueue_output_ready = ~writeResponseQueue_empty & io_coordinator_writeResponse_valid; // @[ExternalMemoryInterface.scala 224:37 263:37]
  always @(posedge clock) begin
    if (reset) begin // @[ExternalMemoryInterface.scala 116:27]
      readQueued <= 1'h0; // @[ExternalMemoryInterface.scala 116:27]
    end else if (~readQueue_full) begin // @[ExternalMemoryInterface.scala 118:25]
      if (instructionOrReadDataQueue_output_valid) begin // @[ExternalMemoryInterface.scala 119:33]
        if (io_coordinator_readAddress_ready) begin // @[ExternalMemoryInterface.scala 136:46]
          readQueued <= 1'h0; // @[ExternalMemoryInterface.scala 138:20]
        end else begin
          readQueued <= 1'h1; // @[ExternalMemoryInterface.scala 135:18]
        end
      end
    end
    if (reset) begin // @[ExternalMemoryInterface.scala 117:25]
      burstLen <= 8'h0; // @[ExternalMemoryInterface.scala 117:25]
    end else if (~readQueue_full) begin // @[ExternalMemoryInterface.scala 118:25]
      if (~readQueue_empty) begin // @[ExternalMemoryInterface.scala 141:28]
        if (io_coordinator_read_valid) begin // @[ExternalMemoryInterface.scala 147:39]
          burstLen <= _GEN_20;
        end
      end
    end
    if (reset) begin // @[ExternalMemoryInterface.scala 229:30]
      writeQueued <= 1'h0; // @[ExternalMemoryInterface.scala 229:30]
    end else if (io_dataWriteRequests_valid) begin // @[ExternalMemoryInterface.scala 230:38]
      if (io_coordinator_writeAddress_ready) begin // @[ExternalMemoryInterface.scala 247:47]
        writeQueued <= 1'h0; // @[ExternalMemoryInterface.scala 249:21]
      end else begin
        writeQueued <= 1'h1; // @[ExternalMemoryInterface.scala 245:21]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  readQueued = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  burstLen = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  writeQueued = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CSRReservationStation(
  input         clock,
  input         reset,
  output        io_decoderInput_0_ready,
  input         io_decoderInput_0_valid,
  input         io_decoderInput_0_bits_sourceTag_threadId,
  input  [3:0]  io_decoderInput_0_bits_sourceTag_id,
  input         io_decoderInput_0_bits_destinationTag_threadId,
  input  [3:0]  io_decoderInput_0_bits_destinationTag_id,
  input  [63:0] io_decoderInput_0_bits_value,
  input         io_decoderInput_0_bits_ready,
  input  [11:0] io_decoderInput_0_bits_address,
  input  [1:0]  io_decoderInput_0_bits_csrAccessType,
  input         io_toCSR_ready,
  output        io_toCSR_valid,
  output [11:0] io_toCSR_bits_address,
  output [63:0] io_toCSR_bits_value,
  output        io_toCSR_bits_destinationTag_threadId,
  output [3:0]  io_toCSR_bits_destinationTag_id,
  output [1:0]  io_toCSR_bits_csrAccessType,
  input         io_output_outputs_valid,
  input  [63:0] io_output_outputs_bits_value,
  input         io_output_outputs_bits_tag_threadId,
  input  [3:0]  io_output_outputs_bits_tag_id,
  output        io_empty
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] head; // @[CSRReservationStation.scala 30:29]
  reg [1:0] tail; // @[CSRReservationStation.scala 31:29]
  reg  buf_0_valid; // @[CSRReservationStation.scala 32:28]
  reg  buf_0_sourceTag_threadId; // @[CSRReservationStation.scala 32:28]
  reg [3:0] buf_0_sourceTag_id; // @[CSRReservationStation.scala 32:28]
  reg [63:0] buf_0_value; // @[CSRReservationStation.scala 32:28]
  reg  buf_0_ready; // @[CSRReservationStation.scala 32:28]
  reg  buf_0_destinationTag_threadId; // @[CSRReservationStation.scala 32:28]
  reg [3:0] buf_0_destinationTag_id; // @[CSRReservationStation.scala 32:28]
  reg [11:0] buf_0_address; // @[CSRReservationStation.scala 32:28]
  reg [1:0] buf_0_csrAccessType; // @[CSRReservationStation.scala 32:28]
  reg  buf_1_valid; // @[CSRReservationStation.scala 32:28]
  reg  buf_1_sourceTag_threadId; // @[CSRReservationStation.scala 32:28]
  reg [3:0] buf_1_sourceTag_id; // @[CSRReservationStation.scala 32:28]
  reg [63:0] buf_1_value; // @[CSRReservationStation.scala 32:28]
  reg  buf_1_ready; // @[CSRReservationStation.scala 32:28]
  reg  buf_1_destinationTag_threadId; // @[CSRReservationStation.scala 32:28]
  reg [3:0] buf_1_destinationTag_id; // @[CSRReservationStation.scala 32:28]
  reg [11:0] buf_1_address; // @[CSRReservationStation.scala 32:28]
  reg [1:0] buf_1_csrAccessType; // @[CSRReservationStation.scala 32:28]
  reg  buf_2_valid; // @[CSRReservationStation.scala 32:28]
  reg  buf_2_sourceTag_threadId; // @[CSRReservationStation.scala 32:28]
  reg [3:0] buf_2_sourceTag_id; // @[CSRReservationStation.scala 32:28]
  reg [63:0] buf_2_value; // @[CSRReservationStation.scala 32:28]
  reg  buf_2_ready; // @[CSRReservationStation.scala 32:28]
  reg  buf_2_destinationTag_threadId; // @[CSRReservationStation.scala 32:28]
  reg [3:0] buf_2_destinationTag_id; // @[CSRReservationStation.scala 32:28]
  reg [11:0] buf_2_address; // @[CSRReservationStation.scala 32:28]
  reg [1:0] buf_2_csrAccessType; // @[CSRReservationStation.scala 32:28]
  reg  buf_3_valid; // @[CSRReservationStation.scala 32:28]
  reg  buf_3_sourceTag_threadId; // @[CSRReservationStation.scala 32:28]
  reg [3:0] buf_3_sourceTag_id; // @[CSRReservationStation.scala 32:28]
  reg [63:0] buf_3_value; // @[CSRReservationStation.scala 32:28]
  reg  buf_3_ready; // @[CSRReservationStation.scala 32:28]
  reg  buf_3_destinationTag_threadId; // @[CSRReservationStation.scala 32:28]
  reg [3:0] buf_3_destinationTag_id; // @[CSRReservationStation.scala 32:28]
  reg [11:0] buf_3_address; // @[CSRReservationStation.scala 32:28]
  reg [1:0] buf_3_csrAccessType; // @[CSRReservationStation.scala 32:28]
  wire [1:0] _io_decoderInput_0_ready_T_1 = head + 2'h1; // @[CSRReservationStation.scala 39:37]
  wire  _T = io_decoderInput_0_ready & io_decoderInput_0_valid; // @[CSRReservationStation.scala 40:18]
  wire  _GEN_0 = 2'h0 == head | buf_0_valid; // @[CSRReservationStation.scala 41:{24,24} 32:28]
  wire  _GEN_1 = 2'h1 == head | buf_1_valid; // @[CSRReservationStation.scala 41:{24,24} 32:28]
  wire  _GEN_2 = 2'h2 == head | buf_2_valid; // @[CSRReservationStation.scala 41:{24,24} 32:28]
  wire  _GEN_3 = 2'h3 == head | buf_3_valid; // @[CSRReservationStation.scala 41:{24,24} 32:28]
  wire [63:0] _GEN_12 = 2'h0 == head ? io_decoderInput_0_bits_value : buf_0_value; // @[CSRReservationStation.scala 41:{24,24} 32:28]
  wire [63:0] _GEN_13 = 2'h1 == head ? io_decoderInput_0_bits_value : buf_1_value; // @[CSRReservationStation.scala 41:{24,24} 32:28]
  wire [63:0] _GEN_14 = 2'h2 == head ? io_decoderInput_0_bits_value : buf_2_value; // @[CSRReservationStation.scala 41:{24,24} 32:28]
  wire [63:0] _GEN_15 = 2'h3 == head ? io_decoderInput_0_bits_value : buf_3_value; // @[CSRReservationStation.scala 41:{24,24} 32:28]
  wire  _GEN_16 = 2'h0 == head ? io_decoderInput_0_bits_ready : buf_0_ready; // @[CSRReservationStation.scala 41:{24,24} 32:28]
  wire  _GEN_17 = 2'h1 == head ? io_decoderInput_0_bits_ready : buf_1_ready; // @[CSRReservationStation.scala 41:{24,24} 32:28]
  wire  _GEN_18 = 2'h2 == head ? io_decoderInput_0_bits_ready : buf_2_ready; // @[CSRReservationStation.scala 41:{24,24} 32:28]
  wire  _GEN_19 = 2'h3 == head ? io_decoderInput_0_bits_ready : buf_3_ready; // @[CSRReservationStation.scala 41:{24,24} 32:28]
  wire  _GEN_36 = io_decoderInput_0_ready & io_decoderInput_0_valid ? _GEN_0 : buf_0_valid; // @[CSRReservationStation.scala 32:28 40:30]
  wire  _GEN_37 = io_decoderInput_0_ready & io_decoderInput_0_valid ? _GEN_1 : buf_1_valid; // @[CSRReservationStation.scala 32:28 40:30]
  wire  _GEN_38 = io_decoderInput_0_ready & io_decoderInput_0_valid ? _GEN_2 : buf_2_valid; // @[CSRReservationStation.scala 32:28 40:30]
  wire  _GEN_39 = io_decoderInput_0_ready & io_decoderInput_0_valid ? _GEN_3 : buf_3_valid; // @[CSRReservationStation.scala 32:28 40:30]
  wire [63:0] _GEN_48 = io_decoderInput_0_ready & io_decoderInput_0_valid ? _GEN_12 : buf_0_value; // @[CSRReservationStation.scala 32:28 40:30]
  wire [63:0] _GEN_49 = io_decoderInput_0_ready & io_decoderInput_0_valid ? _GEN_13 : buf_1_value; // @[CSRReservationStation.scala 32:28 40:30]
  wire [63:0] _GEN_50 = io_decoderInput_0_ready & io_decoderInput_0_valid ? _GEN_14 : buf_2_value; // @[CSRReservationStation.scala 32:28 40:30]
  wire [63:0] _GEN_51 = io_decoderInput_0_ready & io_decoderInput_0_valid ? _GEN_15 : buf_3_value; // @[CSRReservationStation.scala 32:28 40:30]
  wire  _GEN_52 = io_decoderInput_0_ready & io_decoderInput_0_valid ? _GEN_16 : buf_0_ready; // @[CSRReservationStation.scala 32:28 40:30]
  wire  _GEN_53 = io_decoderInput_0_ready & io_decoderInput_0_valid ? _GEN_17 : buf_1_ready; // @[CSRReservationStation.scala 32:28 40:30]
  wire  _GEN_54 = io_decoderInput_0_ready & io_decoderInput_0_valid ? _GEN_18 : buf_2_ready; // @[CSRReservationStation.scala 32:28 40:30]
  wire  _GEN_55 = io_decoderInput_0_ready & io_decoderInput_0_valid ? _GEN_19 : buf_3_ready; // @[CSRReservationStation.scala 32:28 40:30]
  wire  _GEN_73 = 2'h1 == tail ? buf_1_ready : buf_0_ready; // @[CSRReservationStation.scala 57:{22,22}]
  wire  _GEN_74 = 2'h2 == tail ? buf_2_ready : _GEN_73; // @[CSRReservationStation.scala 57:{22,22}]
  wire  _GEN_75 = 2'h3 == tail ? buf_3_ready : _GEN_74; // @[CSRReservationStation.scala 57:{22,22}]
  wire [63:0] _GEN_77 = 2'h1 == tail ? buf_1_value : buf_0_value; // @[CSRReservationStation.scala 59:{25,25}]
  wire [63:0] _GEN_78 = 2'h2 == tail ? buf_2_value : _GEN_77; // @[CSRReservationStation.scala 59:{25,25}]
  wire [11:0] _GEN_81 = 2'h1 == tail ? buf_1_address : buf_0_address; // @[CSRReservationStation.scala 60:{27,27}]
  wire [11:0] _GEN_82 = 2'h2 == tail ? buf_2_address : _GEN_81; // @[CSRReservationStation.scala 60:{27,27}]
  wire  _GEN_85 = 2'h1 == tail ? buf_1_destinationTag_threadId : buf_0_destinationTag_threadId; // @[CSRReservationStation.scala 61:{34,34}]
  wire  _GEN_86 = 2'h2 == tail ? buf_2_destinationTag_threadId : _GEN_85; // @[CSRReservationStation.scala 61:{34,34}]
  wire [3:0] _GEN_89 = 2'h1 == tail ? buf_1_destinationTag_id : buf_0_destinationTag_id; // @[CSRReservationStation.scala 61:{34,34}]
  wire [3:0] _GEN_90 = 2'h2 == tail ? buf_2_destinationTag_id : _GEN_89; // @[CSRReservationStation.scala 61:{34,34}]
  wire [1:0] _GEN_93 = 2'h1 == tail ? buf_1_csrAccessType : buf_0_csrAccessType; // @[CSRReservationStation.scala 62:{33,33}]
  wire [1:0] _GEN_94 = 2'h2 == tail ? buf_2_csrAccessType : _GEN_93; // @[CSRReservationStation.scala 62:{33,33}]
  wire [1:0] _tail_T_1 = tail + 2'h1; // @[CSRReservationStation.scala 64:20]
  wire  _T_10 = buf_0_sourceTag_id == io_output_outputs_bits_tag_id & buf_0_sourceTag_threadId ==
    io_output_outputs_bits_tag_threadId; // @[Tag.scala 13:25]
  wire  _GEN_117 = buf_0_valid & ~buf_0_ready & _T_10 | _GEN_52; // @[CSRReservationStation.scala 71:79 73:17]
  wire  _T_16 = buf_1_sourceTag_id == io_output_outputs_bits_tag_id & buf_1_sourceTag_threadId ==
    io_output_outputs_bits_tag_threadId; // @[Tag.scala 13:25]
  wire  _GEN_119 = buf_1_valid & ~buf_1_ready & _T_16 | _GEN_53; // @[CSRReservationStation.scala 71:79 73:17]
  wire  _T_22 = buf_2_sourceTag_id == io_output_outputs_bits_tag_id & buf_2_sourceTag_threadId ==
    io_output_outputs_bits_tag_threadId; // @[Tag.scala 13:25]
  wire  _GEN_121 = buf_2_valid & ~buf_2_ready & _T_22 | _GEN_54; // @[CSRReservationStation.scala 71:79 73:17]
  wire  _T_28 = buf_3_sourceTag_id == io_output_outputs_bits_tag_id & buf_3_sourceTag_threadId ==
    io_output_outputs_bits_tag_threadId; // @[Tag.scala 13:25]
  wire  _GEN_123 = buf_3_valid & ~buf_3_ready & _T_28 | _GEN_55; // @[CSRReservationStation.scala 71:79 73:17]
  assign io_decoderInput_0_ready = tail != _io_decoderInput_0_ready_T_1; // @[CSRReservationStation.scala 39:21]
  assign io_toCSR_valid = tail != head & _GEN_75; // @[CSRReservationStation.scala 57:22]
  assign io_toCSR_bits_address = 2'h3 == tail ? buf_3_address : _GEN_82; // @[CSRReservationStation.scala 60:{27,27}]
  assign io_toCSR_bits_value = 2'h3 == tail ? buf_3_value : _GEN_78; // @[CSRReservationStation.scala 59:{25,25}]
  assign io_toCSR_bits_destinationTag_threadId = 2'h3 == tail ? buf_3_destinationTag_threadId : _GEN_86; // @[CSRReservationStation.scala 61:{34,34}]
  assign io_toCSR_bits_destinationTag_id = 2'h3 == tail ? buf_3_destinationTag_id : _GEN_90; // @[CSRReservationStation.scala 61:{34,34}]
  assign io_toCSR_bits_csrAccessType = 2'h3 == tail ? buf_3_csrAccessType : _GEN_94; // @[CSRReservationStation.scala 62:{33,33}]
  assign io_empty = head == tail; // @[CSRReservationStation.scala 35:20]
  always @(posedge clock) begin
    if (reset) begin // @[CSRReservationStation.scala 30:29]
      head <= 2'h0; // @[CSRReservationStation.scala 30:29]
    end else if (_T) begin // @[CSRReservationStation.scala 53:22]
      head <= _io_decoderInput_0_ready_T_1;
    end
    if (reset) begin // @[CSRReservationStation.scala 31:29]
      tail <= 2'h0; // @[CSRReservationStation.scala 31:29]
    end else if (tail != head & _GEN_75) begin // @[CSRReservationStation.scala 57:42]
      if (io_toCSR_ready) begin // @[CSRReservationStation.scala 63:26]
        tail <= _tail_T_1; // @[CSRReservationStation.scala 64:12]
      end
    end
    if (reset) begin // @[CSRReservationStation.scala 32:28]
      buf_0_valid <= 1'h0; // @[CSRReservationStation.scala 32:28]
    end else if (tail != head & _GEN_75) begin // @[CSRReservationStation.scala 57:42]
      if (io_toCSR_ready) begin // @[CSRReservationStation.scala 63:26]
        if (2'h0 == tail) begin // @[CSRReservationStation.scala 65:23]
          buf_0_valid <= 1'h0; // @[CSRReservationStation.scala 65:23]
        end else begin
          buf_0_valid <= _GEN_36;
        end
      end else begin
        buf_0_valid <= _GEN_36;
      end
    end else begin
      buf_0_valid <= _GEN_36;
    end
    if (io_decoderInput_0_ready & io_decoderInput_0_valid) begin // @[CSRReservationStation.scala 40:30]
      if (2'h0 == head) begin // @[CSRReservationStation.scala 41:24]
        buf_0_sourceTag_threadId <= io_decoderInput_0_bits_sourceTag_threadId; // @[CSRReservationStation.scala 41:24]
      end
    end
    if (io_decoderInput_0_ready & io_decoderInput_0_valid) begin // @[CSRReservationStation.scala 40:30]
      if (2'h0 == head) begin // @[CSRReservationStation.scala 41:24]
        buf_0_sourceTag_id <= io_decoderInput_0_bits_sourceTag_id; // @[CSRReservationStation.scala 41:24]
      end
    end
    if (io_output_outputs_valid) begin // @[CSRReservationStation.scala 69:33]
      if (buf_0_valid & ~buf_0_ready & _T_10) begin // @[CSRReservationStation.scala 71:79]
        buf_0_value <= io_output_outputs_bits_value; // @[CSRReservationStation.scala 72:17]
      end else begin
        buf_0_value <= _GEN_48;
      end
    end else begin
      buf_0_value <= _GEN_48;
    end
    if (io_output_outputs_valid) begin // @[CSRReservationStation.scala 69:33]
      buf_0_ready <= _GEN_117;
    end else if (io_decoderInput_0_ready & io_decoderInput_0_valid) begin // @[CSRReservationStation.scala 40:30]
      if (2'h0 == head) begin // @[CSRReservationStation.scala 41:24]
        buf_0_ready <= io_decoderInput_0_bits_ready; // @[CSRReservationStation.scala 41:24]
      end
    end
    if (io_decoderInput_0_ready & io_decoderInput_0_valid) begin // @[CSRReservationStation.scala 40:30]
      if (2'h0 == head) begin // @[CSRReservationStation.scala 41:24]
        buf_0_destinationTag_threadId <= io_decoderInput_0_bits_destinationTag_threadId; // @[CSRReservationStation.scala 41:24]
      end
    end
    if (io_decoderInput_0_ready & io_decoderInput_0_valid) begin // @[CSRReservationStation.scala 40:30]
      if (2'h0 == head) begin // @[CSRReservationStation.scala 41:24]
        buf_0_destinationTag_id <= io_decoderInput_0_bits_destinationTag_id; // @[CSRReservationStation.scala 41:24]
      end
    end
    if (io_decoderInput_0_ready & io_decoderInput_0_valid) begin // @[CSRReservationStation.scala 40:30]
      if (2'h0 == head) begin // @[CSRReservationStation.scala 41:24]
        buf_0_address <= io_decoderInput_0_bits_address; // @[CSRReservationStation.scala 41:24]
      end
    end
    if (io_decoderInput_0_ready & io_decoderInput_0_valid) begin // @[CSRReservationStation.scala 40:30]
      if (2'h0 == head) begin // @[CSRReservationStation.scala 41:24]
        buf_0_csrAccessType <= io_decoderInput_0_bits_csrAccessType; // @[CSRReservationStation.scala 41:24]
      end
    end
    if (reset) begin // @[CSRReservationStation.scala 32:28]
      buf_1_valid <= 1'h0; // @[CSRReservationStation.scala 32:28]
    end else if (tail != head & _GEN_75) begin // @[CSRReservationStation.scala 57:42]
      if (io_toCSR_ready) begin // @[CSRReservationStation.scala 63:26]
        if (2'h1 == tail) begin // @[CSRReservationStation.scala 65:23]
          buf_1_valid <= 1'h0; // @[CSRReservationStation.scala 65:23]
        end else begin
          buf_1_valid <= _GEN_37;
        end
      end else begin
        buf_1_valid <= _GEN_37;
      end
    end else begin
      buf_1_valid <= _GEN_37;
    end
    if (io_decoderInput_0_ready & io_decoderInput_0_valid) begin // @[CSRReservationStation.scala 40:30]
      if (2'h1 == head) begin // @[CSRReservationStation.scala 41:24]
        buf_1_sourceTag_threadId <= io_decoderInput_0_bits_sourceTag_threadId; // @[CSRReservationStation.scala 41:24]
      end
    end
    if (io_decoderInput_0_ready & io_decoderInput_0_valid) begin // @[CSRReservationStation.scala 40:30]
      if (2'h1 == head) begin // @[CSRReservationStation.scala 41:24]
        buf_1_sourceTag_id <= io_decoderInput_0_bits_sourceTag_id; // @[CSRReservationStation.scala 41:24]
      end
    end
    if (io_output_outputs_valid) begin // @[CSRReservationStation.scala 69:33]
      if (buf_1_valid & ~buf_1_ready & _T_16) begin // @[CSRReservationStation.scala 71:79]
        buf_1_value <= io_output_outputs_bits_value; // @[CSRReservationStation.scala 72:17]
      end else begin
        buf_1_value <= _GEN_49;
      end
    end else begin
      buf_1_value <= _GEN_49;
    end
    if (io_output_outputs_valid) begin // @[CSRReservationStation.scala 69:33]
      buf_1_ready <= _GEN_119;
    end else if (io_decoderInput_0_ready & io_decoderInput_0_valid) begin // @[CSRReservationStation.scala 40:30]
      if (2'h1 == head) begin // @[CSRReservationStation.scala 41:24]
        buf_1_ready <= io_decoderInput_0_bits_ready; // @[CSRReservationStation.scala 41:24]
      end
    end
    if (io_decoderInput_0_ready & io_decoderInput_0_valid) begin // @[CSRReservationStation.scala 40:30]
      if (2'h1 == head) begin // @[CSRReservationStation.scala 41:24]
        buf_1_destinationTag_threadId <= io_decoderInput_0_bits_destinationTag_threadId; // @[CSRReservationStation.scala 41:24]
      end
    end
    if (io_decoderInput_0_ready & io_decoderInput_0_valid) begin // @[CSRReservationStation.scala 40:30]
      if (2'h1 == head) begin // @[CSRReservationStation.scala 41:24]
        buf_1_destinationTag_id <= io_decoderInput_0_bits_destinationTag_id; // @[CSRReservationStation.scala 41:24]
      end
    end
    if (io_decoderInput_0_ready & io_decoderInput_0_valid) begin // @[CSRReservationStation.scala 40:30]
      if (2'h1 == head) begin // @[CSRReservationStation.scala 41:24]
        buf_1_address <= io_decoderInput_0_bits_address; // @[CSRReservationStation.scala 41:24]
      end
    end
    if (io_decoderInput_0_ready & io_decoderInput_0_valid) begin // @[CSRReservationStation.scala 40:30]
      if (2'h1 == head) begin // @[CSRReservationStation.scala 41:24]
        buf_1_csrAccessType <= io_decoderInput_0_bits_csrAccessType; // @[CSRReservationStation.scala 41:24]
      end
    end
    if (reset) begin // @[CSRReservationStation.scala 32:28]
      buf_2_valid <= 1'h0; // @[CSRReservationStation.scala 32:28]
    end else if (tail != head & _GEN_75) begin // @[CSRReservationStation.scala 57:42]
      if (io_toCSR_ready) begin // @[CSRReservationStation.scala 63:26]
        if (2'h2 == tail) begin // @[CSRReservationStation.scala 65:23]
          buf_2_valid <= 1'h0; // @[CSRReservationStation.scala 65:23]
        end else begin
          buf_2_valid <= _GEN_38;
        end
      end else begin
        buf_2_valid <= _GEN_38;
      end
    end else begin
      buf_2_valid <= _GEN_38;
    end
    if (io_decoderInput_0_ready & io_decoderInput_0_valid) begin // @[CSRReservationStation.scala 40:30]
      if (2'h2 == head) begin // @[CSRReservationStation.scala 41:24]
        buf_2_sourceTag_threadId <= io_decoderInput_0_bits_sourceTag_threadId; // @[CSRReservationStation.scala 41:24]
      end
    end
    if (io_decoderInput_0_ready & io_decoderInput_0_valid) begin // @[CSRReservationStation.scala 40:30]
      if (2'h2 == head) begin // @[CSRReservationStation.scala 41:24]
        buf_2_sourceTag_id <= io_decoderInput_0_bits_sourceTag_id; // @[CSRReservationStation.scala 41:24]
      end
    end
    if (io_output_outputs_valid) begin // @[CSRReservationStation.scala 69:33]
      if (buf_2_valid & ~buf_2_ready & _T_22) begin // @[CSRReservationStation.scala 71:79]
        buf_2_value <= io_output_outputs_bits_value; // @[CSRReservationStation.scala 72:17]
      end else begin
        buf_2_value <= _GEN_50;
      end
    end else begin
      buf_2_value <= _GEN_50;
    end
    if (io_output_outputs_valid) begin // @[CSRReservationStation.scala 69:33]
      buf_2_ready <= _GEN_121;
    end else if (io_decoderInput_0_ready & io_decoderInput_0_valid) begin // @[CSRReservationStation.scala 40:30]
      if (2'h2 == head) begin // @[CSRReservationStation.scala 41:24]
        buf_2_ready <= io_decoderInput_0_bits_ready; // @[CSRReservationStation.scala 41:24]
      end
    end
    if (io_decoderInput_0_ready & io_decoderInput_0_valid) begin // @[CSRReservationStation.scala 40:30]
      if (2'h2 == head) begin // @[CSRReservationStation.scala 41:24]
        buf_2_destinationTag_threadId <= io_decoderInput_0_bits_destinationTag_threadId; // @[CSRReservationStation.scala 41:24]
      end
    end
    if (io_decoderInput_0_ready & io_decoderInput_0_valid) begin // @[CSRReservationStation.scala 40:30]
      if (2'h2 == head) begin // @[CSRReservationStation.scala 41:24]
        buf_2_destinationTag_id <= io_decoderInput_0_bits_destinationTag_id; // @[CSRReservationStation.scala 41:24]
      end
    end
    if (io_decoderInput_0_ready & io_decoderInput_0_valid) begin // @[CSRReservationStation.scala 40:30]
      if (2'h2 == head) begin // @[CSRReservationStation.scala 41:24]
        buf_2_address <= io_decoderInput_0_bits_address; // @[CSRReservationStation.scala 41:24]
      end
    end
    if (io_decoderInput_0_ready & io_decoderInput_0_valid) begin // @[CSRReservationStation.scala 40:30]
      if (2'h2 == head) begin // @[CSRReservationStation.scala 41:24]
        buf_2_csrAccessType <= io_decoderInput_0_bits_csrAccessType; // @[CSRReservationStation.scala 41:24]
      end
    end
    if (reset) begin // @[CSRReservationStation.scala 32:28]
      buf_3_valid <= 1'h0; // @[CSRReservationStation.scala 32:28]
    end else if (tail != head & _GEN_75) begin // @[CSRReservationStation.scala 57:42]
      if (io_toCSR_ready) begin // @[CSRReservationStation.scala 63:26]
        if (2'h3 == tail) begin // @[CSRReservationStation.scala 65:23]
          buf_3_valid <= 1'h0; // @[CSRReservationStation.scala 65:23]
        end else begin
          buf_3_valid <= _GEN_39;
        end
      end else begin
        buf_3_valid <= _GEN_39;
      end
    end else begin
      buf_3_valid <= _GEN_39;
    end
    if (io_decoderInput_0_ready & io_decoderInput_0_valid) begin // @[CSRReservationStation.scala 40:30]
      if (2'h3 == head) begin // @[CSRReservationStation.scala 41:24]
        buf_3_sourceTag_threadId <= io_decoderInput_0_bits_sourceTag_threadId; // @[CSRReservationStation.scala 41:24]
      end
    end
    if (io_decoderInput_0_ready & io_decoderInput_0_valid) begin // @[CSRReservationStation.scala 40:30]
      if (2'h3 == head) begin // @[CSRReservationStation.scala 41:24]
        buf_3_sourceTag_id <= io_decoderInput_0_bits_sourceTag_id; // @[CSRReservationStation.scala 41:24]
      end
    end
    if (io_output_outputs_valid) begin // @[CSRReservationStation.scala 69:33]
      if (buf_3_valid & ~buf_3_ready & _T_28) begin // @[CSRReservationStation.scala 71:79]
        buf_3_value <= io_output_outputs_bits_value; // @[CSRReservationStation.scala 72:17]
      end else begin
        buf_3_value <= _GEN_51;
      end
    end else begin
      buf_3_value <= _GEN_51;
    end
    if (io_output_outputs_valid) begin // @[CSRReservationStation.scala 69:33]
      buf_3_ready <= _GEN_123;
    end else if (io_decoderInput_0_ready & io_decoderInput_0_valid) begin // @[CSRReservationStation.scala 40:30]
      if (2'h3 == head) begin // @[CSRReservationStation.scala 41:24]
        buf_3_ready <= io_decoderInput_0_bits_ready; // @[CSRReservationStation.scala 41:24]
      end
    end
    if (io_decoderInput_0_ready & io_decoderInput_0_valid) begin // @[CSRReservationStation.scala 40:30]
      if (2'h3 == head) begin // @[CSRReservationStation.scala 41:24]
        buf_3_destinationTag_threadId <= io_decoderInput_0_bits_destinationTag_threadId; // @[CSRReservationStation.scala 41:24]
      end
    end
    if (io_decoderInput_0_ready & io_decoderInput_0_valid) begin // @[CSRReservationStation.scala 40:30]
      if (2'h3 == head) begin // @[CSRReservationStation.scala 41:24]
        buf_3_destinationTag_id <= io_decoderInput_0_bits_destinationTag_id; // @[CSRReservationStation.scala 41:24]
      end
    end
    if (io_decoderInput_0_ready & io_decoderInput_0_valid) begin // @[CSRReservationStation.scala 40:30]
      if (2'h3 == head) begin // @[CSRReservationStation.scala 41:24]
        buf_3_address <= io_decoderInput_0_bits_address; // @[CSRReservationStation.scala 41:24]
      end
    end
    if (io_decoderInput_0_ready & io_decoderInput_0_valid) begin // @[CSRReservationStation.scala 40:30]
      if (2'h3 == head) begin // @[CSRReservationStation.scala 41:24]
        buf_3_csrAccessType <= io_decoderInput_0_bits_csrAccessType; // @[CSRReservationStation.scala 41:24]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  head = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  tail = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  buf_0_valid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  buf_0_sourceTag_threadId = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  buf_0_sourceTag_id = _RAND_4[3:0];
  _RAND_5 = {2{`RANDOM}};
  buf_0_value = _RAND_5[63:0];
  _RAND_6 = {1{`RANDOM}};
  buf_0_ready = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  buf_0_destinationTag_threadId = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  buf_0_destinationTag_id = _RAND_8[3:0];
  _RAND_9 = {1{`RANDOM}};
  buf_0_address = _RAND_9[11:0];
  _RAND_10 = {1{`RANDOM}};
  buf_0_csrAccessType = _RAND_10[1:0];
  _RAND_11 = {1{`RANDOM}};
  buf_1_valid = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  buf_1_sourceTag_threadId = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  buf_1_sourceTag_id = _RAND_13[3:0];
  _RAND_14 = {2{`RANDOM}};
  buf_1_value = _RAND_14[63:0];
  _RAND_15 = {1{`RANDOM}};
  buf_1_ready = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  buf_1_destinationTag_threadId = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  buf_1_destinationTag_id = _RAND_17[3:0];
  _RAND_18 = {1{`RANDOM}};
  buf_1_address = _RAND_18[11:0];
  _RAND_19 = {1{`RANDOM}};
  buf_1_csrAccessType = _RAND_19[1:0];
  _RAND_20 = {1{`RANDOM}};
  buf_2_valid = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  buf_2_sourceTag_threadId = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  buf_2_sourceTag_id = _RAND_22[3:0];
  _RAND_23 = {2{`RANDOM}};
  buf_2_value = _RAND_23[63:0];
  _RAND_24 = {1{`RANDOM}};
  buf_2_ready = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  buf_2_destinationTag_threadId = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  buf_2_destinationTag_id = _RAND_26[3:0];
  _RAND_27 = {1{`RANDOM}};
  buf_2_address = _RAND_27[11:0];
  _RAND_28 = {1{`RANDOM}};
  buf_2_csrAccessType = _RAND_28[1:0];
  _RAND_29 = {1{`RANDOM}};
  buf_3_valid = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  buf_3_sourceTag_threadId = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  buf_3_sourceTag_id = _RAND_31[3:0];
  _RAND_32 = {2{`RANDOM}};
  buf_3_value = _RAND_32[63:0];
  _RAND_33 = {1{`RANDOM}};
  buf_3_ready = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  buf_3_destinationTag_threadId = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  buf_3_destinationTag_id = _RAND_35[3:0];
  _RAND_36 = {1{`RANDOM}};
  buf_3_address = _RAND_36[11:0];
  _RAND_37 = {1{`RANDOM}};
  buf_3_csrAccessType = _RAND_37[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RetireCounter(
  input         clock,
  input         reset,
  input  [1:0]  io_retireInCycle,
  output [63:0] io_count
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] c; // @[RetireCounter.scala 14:18]
  wire [63:0] _GEN_0 = {{62'd0}, io_retireInCycle}; // @[RetireCounter.scala 15:10]
  wire [63:0] _c_T_1 = c + _GEN_0; // @[RetireCounter.scala 15:10]
  assign io_count = c; // @[RetireCounter.scala 16:12]
  always @(posedge clock) begin
    if (reset) begin // @[RetireCounter.scala 14:18]
      c <= 64'h0; // @[RetireCounter.scala 14:18]
    end else begin
      c <= _c_T_1; // @[RetireCounter.scala 15:5]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  c = _RAND_0[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CycleCounter(
  input         clock,
  input         reset,
  output [63:0] count
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] c; // @[CycleCounter.scala 8:26]
  wire [63:0] _c_T_1 = c + 64'h1; // @[CycleCounter.scala 9:10]
  assign count = c; // @[CycleCounter.scala 10:9]
  always @(posedge clock) begin
    if (reset) begin // @[CycleCounter.scala 8:26]
      c <= 64'h0; // @[CycleCounter.scala 8:26]
    end else begin
      c <= _c_T_1; // @[CycleCounter.scala 9:5]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  c = _RAND_0[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CSR(
  input         clock,
  input         reset,
  output        io_decoderInput_ready,
  input         io_decoderInput_valid,
  input  [11:0] io_decoderInput_bits_address,
  input  [63:0] io_decoderInput_bits_value,
  input         io_decoderInput_bits_destinationTag_threadId,
  input  [3:0]  io_decoderInput_bits_destinationTag_id,
  input  [1:0]  io_decoderInput_bits_csrAccessType,
  input         io_CSROutput_ready,
  output        io_CSROutput_valid,
  output [63:0] io_CSROutput_bits_value,
  output        io_CSROutput_bits_isError,
  output        io_CSROutput_bits_tag_threadId,
  output [3:0]  io_CSROutput_bits_tag_id,
  output [63:0] io_fetch_mtvec,
  output [63:0] io_fetch_mepc,
  output [63:0] io_fetch_mcause,
  input  [1:0]  io_reorderBuffer_retireCount
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  retireCounter_clock; // @[CSR.scala 32:29]
  wire  retireCounter_reset; // @[CSR.scala 32:29]
  wire [1:0] retireCounter_io_retireInCycle; // @[CSR.scala 32:29]
  wire [63:0] retireCounter_io_count; // @[CSR.scala 32:29]
  wire  cycleCounter_clock; // @[CSR.scala 34:28]
  wire  cycleCounter_reset; // @[CSR.scala 34:28]
  wire [63:0] cycleCounter_count; // @[CSR.scala 34:28]
  reg [63:0] mtvec; // @[CSR.scala 36:22]
  reg [63:0] mepc; // @[CSR.scala 38:21]
  reg [63:0] mcause; // @[CSR.scala 40:23]
  reg [63:0] mstatus; // @[CSR.scala 42:24]
  wire  _T_8 = io_CSROutput_ready & io_CSROutput_valid; // @[CSR.scala 56:31]
  wire [63:0] _mtvec_T_3 = mtvec | io_decoderInput_bits_value; // @[CSR.scala 62:52]
  wire [63:0] _mtvec_T_5 = mtvec & io_decoderInput_bits_value; // @[CSR.scala 63:54]
  wire [63:0] _mtvec_T_7 = 2'h0 == io_decoderInput_bits_csrAccessType ? io_decoderInput_bits_value : 64'h0; // @[Mux.scala 81:58]
  wire [63:0] _mtvec_T_9 = 2'h1 == io_decoderInput_bits_csrAccessType ? _mtvec_T_3 : _mtvec_T_7; // @[Mux.scala 81:58]
  wire [63:0] _mtvec_T_11 = 2'h2 == io_decoderInput_bits_csrAccessType ? _mtvec_T_5 : _mtvec_T_9; // @[Mux.scala 81:58]
  wire [63:0] _GEN_0 = io_CSROutput_ready & io_CSROutput_valid ? _mtvec_T_11 : mtvec; // @[CSR.scala 56:54 57:15 36:22]
  wire [63:0] _mepc_T_3 = mepc | io_decoderInput_bits_value; // @[CSR.scala 75:51]
  wire [63:0] _mepc_T_5 = mepc & io_decoderInput_bits_value; // @[CSR.scala 76:53]
  wire [63:0] _mepc_T_9 = 2'h1 == io_decoderInput_bits_csrAccessType ? _mepc_T_3 : _mtvec_T_7; // @[Mux.scala 81:58]
  wire [63:0] _mepc_T_11 = 2'h2 == io_decoderInput_bits_csrAccessType ? _mepc_T_5 : _mepc_T_9; // @[Mux.scala 81:58]
  wire [63:0] _GEN_1 = _T_8 ? _mepc_T_11 : mepc; // @[CSR.scala 69:54 70:14 38:21]
  wire [63:0] _mcause_T_3 = mcause | io_decoderInput_bits_value; // @[CSR.scala 88:53]
  wire [63:0] _mcause_T_5 = mcause & io_decoderInput_bits_value; // @[CSR.scala 89:55]
  wire [63:0] _mcause_T_9 = 2'h1 == io_decoderInput_bits_csrAccessType ? _mcause_T_3 : _mtvec_T_7; // @[Mux.scala 81:58]
  wire [63:0] _mcause_T_11 = 2'h2 == io_decoderInput_bits_csrAccessType ? _mcause_T_5 : _mcause_T_9; // @[Mux.scala 81:58]
  wire [63:0] _GEN_2 = _T_8 ? _mcause_T_11 : mcause; // @[CSR.scala 82:54 83:16 40:23]
  wire [63:0] _mstatus_T_3 = mstatus | io_decoderInput_bits_value; // @[CSR.scala 101:54]
  wire [63:0] _mstatus_T_5 = mstatus & io_decoderInput_bits_value; // @[CSR.scala 102:56]
  wire [63:0] _mstatus_T_9 = 2'h1 == io_decoderInput_bits_csrAccessType ? _mstatus_T_3 : _mtvec_T_7; // @[Mux.scala 81:58]
  wire [63:0] _mstatus_T_11 = 2'h2 == io_decoderInput_bits_csrAccessType ? _mstatus_T_5 : _mstatus_T_9; // @[Mux.scala 81:58]
  wire [63:0] _GEN_3 = _T_8 ? _mstatus_T_11 : mstatus; // @[CSR.scala 95:54 96:17 42:24]
  wire [63:0] _GEN_4 = io_decoderInput_bits_address == 12'h300 ? mstatus : 64'h0; // @[CSR.scala 26:27 93:45 94:31]
  wire [63:0] _GEN_5 = io_decoderInput_bits_address == 12'h300 ? _GEN_3 : mstatus; // @[CSR.scala 42:24 93:45]
  wire  _GEN_6 = io_decoderInput_bits_address == 12'h300 ? 1'h0 : 1'h1; // @[CSR.scala 27:29 107:33 93:45]
  wire [63:0] _GEN_7 = io_decoderInput_bits_address == 12'h342 ? mcause : _GEN_4; // @[CSR.scala 80:44 81:31]
  wire [63:0] _GEN_8 = io_decoderInput_bits_address == 12'h342 ? _GEN_2 : mcause; // @[CSR.scala 40:23 80:44]
  wire [63:0] _GEN_9 = io_decoderInput_bits_address == 12'h342 ? mstatus : _GEN_5; // @[CSR.scala 42:24 80:44]
  wire  _GEN_10 = io_decoderInput_bits_address == 12'h342 ? 1'h0 : _GEN_6; // @[CSR.scala 27:29 80:44]
  wire [63:0] _GEN_11 = io_decoderInput_bits_address == 12'h341 ? mepc : _GEN_7; // @[CSR.scala 67:42 68:31]
  wire [63:0] _GEN_12 = io_decoderInput_bits_address == 12'h341 ? _GEN_1 : mepc; // @[CSR.scala 38:21 67:42]
  wire [63:0] _GEN_13 = io_decoderInput_bits_address == 12'h341 ? mcause : _GEN_8; // @[CSR.scala 40:23 67:42]
  wire [63:0] _GEN_14 = io_decoderInput_bits_address == 12'h341 ? mstatus : _GEN_9; // @[CSR.scala 42:24 67:42]
  wire  _GEN_15 = io_decoderInput_bits_address == 12'h341 ? 1'h0 : _GEN_10; // @[CSR.scala 27:29 67:42]
  wire [63:0] _GEN_16 = io_decoderInput_bits_address == 12'h305 ? mtvec : _GEN_11; // @[CSR.scala 54:43 55:31]
  wire [63:0] _GEN_17 = io_decoderInput_bits_address == 12'h305 ? _GEN_0 : mtvec; // @[CSR.scala 36:22 54:43]
  wire [63:0] _GEN_18 = io_decoderInput_bits_address == 12'h305 ? mepc : _GEN_12; // @[CSR.scala 38:21 54:43]
  wire [63:0] _GEN_19 = io_decoderInput_bits_address == 12'h305 ? mcause : _GEN_13; // @[CSR.scala 40:23 54:43]
  wire [63:0] _GEN_20 = io_decoderInput_bits_address == 12'h305 ? mstatus : _GEN_14; // @[CSR.scala 42:24 54:43]
  wire  _GEN_21 = io_decoderInput_bits_address == 12'h305 ? 1'h0 : _GEN_15; // @[CSR.scala 27:29 54:43]
  wire [63:0] _GEN_22 = io_decoderInput_bits_address == 12'hf14 ? 64'h0 : _GEN_16; // @[CSR.scala 52:45 53:31]
  wire [63:0] _GEN_23 = io_decoderInput_bits_address == 12'hf14 ? mtvec : _GEN_17; // @[CSR.scala 36:22 52:45]
  wire [63:0] _GEN_24 = io_decoderInput_bits_address == 12'hf14 ? mepc : _GEN_18; // @[CSR.scala 38:21 52:45]
  wire [63:0] _GEN_25 = io_decoderInput_bits_address == 12'hf14 ? mcause : _GEN_19; // @[CSR.scala 40:23 52:45]
  wire [63:0] _GEN_26 = io_decoderInput_bits_address == 12'hf14 ? mstatus : _GEN_20; // @[CSR.scala 42:24 52:45]
  wire  _GEN_27 = io_decoderInput_bits_address == 12'hf14 ? 1'h0 : _GEN_21; // @[CSR.scala 27:29 52:45]
  wire [63:0] _GEN_28 = io_decoderInput_bits_address == 12'hc02 | io_decoderInput_bits_address == 12'hb02 ?
    retireCounter_io_count : _GEN_22; // @[CSR.scala 50:77 51:31]
  wire  _GEN_33 = io_decoderInput_bits_address == 12'hc02 | io_decoderInput_bits_address == 12'hb02 ? 1'h0 : _GEN_27; // @[CSR.scala 27:29 50:77]
  wire [63:0] _GEN_34 = io_decoderInput_bits_address == 12'hc00 | io_decoderInput_bits_address == 12'hb00 ?
    cycleCounter_count : _GEN_28; // @[CSR.scala 48:67 49:31]
  wire  _GEN_39 = io_decoderInput_bits_address == 12'hc00 | io_decoderInput_bits_address == 12'hb00 ? 1'h0 : _GEN_33; // @[CSR.scala 27:29 48:67]
  RetireCounter retireCounter ( // @[CSR.scala 32:29]
    .clock(retireCounter_clock),
    .reset(retireCounter_reset),
    .io_retireInCycle(retireCounter_io_retireInCycle),
    .io_count(retireCounter_io_count)
  );
  CycleCounter cycleCounter ( // @[CSR.scala 34:28]
    .clock(cycleCounter_clock),
    .reset(cycleCounter_reset),
    .count(cycleCounter_count)
  );
  assign io_decoderInput_ready = io_CSROutput_ready; // @[CSR.scala 23:25]
  assign io_CSROutput_valid = io_decoderInput_valid; // @[CSR.scala 24:22 44:31 46:24]
  assign io_CSROutput_bits_value = io_decoderInput_valid ? _GEN_34 : 64'h0; // @[CSR.scala 26:27 44:31]
  assign io_CSROutput_bits_isError = io_decoderInput_valid & _GEN_39; // @[CSR.scala 27:29 44:31]
  assign io_CSROutput_bits_tag_threadId = io_decoderInput_bits_destinationTag_threadId; // @[CSR.scala 25:25]
  assign io_CSROutput_bits_tag_id = io_decoderInput_bits_destinationTag_id; // @[CSR.scala 25:25]
  assign io_fetch_mtvec = mtvec; // @[CSR.scala 37:18]
  assign io_fetch_mepc = mepc; // @[CSR.scala 39:17]
  assign io_fetch_mcause = mcause; // @[CSR.scala 41:19]
  assign retireCounter_clock = clock;
  assign retireCounter_reset = reset;
  assign retireCounter_io_retireInCycle = io_reorderBuffer_retireCount; // @[CSR.scala 33:34]
  assign cycleCounter_clock = clock;
  assign cycleCounter_reset = reset;
  always @(posedge clock) begin
    if (reset) begin // @[CSR.scala 36:22]
      mtvec <= 64'h0; // @[CSR.scala 36:22]
    end else if (io_decoderInput_valid) begin // @[CSR.scala 44:31]
      if (!(io_decoderInput_bits_address == 12'hc00 | io_decoderInput_bits_address == 12'hb00)) begin // @[CSR.scala 48:67]
        if (!(io_decoderInput_bits_address == 12'hc02 | io_decoderInput_bits_address == 12'hb02)) begin // @[CSR.scala 50:77]
          mtvec <= _GEN_23;
        end
      end
    end
    if (reset) begin // @[CSR.scala 38:21]
      mepc <= 64'h0; // @[CSR.scala 38:21]
    end else if (io_decoderInput_valid) begin // @[CSR.scala 44:31]
      if (!(io_decoderInput_bits_address == 12'hc00 | io_decoderInput_bits_address == 12'hb00)) begin // @[CSR.scala 48:67]
        if (!(io_decoderInput_bits_address == 12'hc02 | io_decoderInput_bits_address == 12'hb02)) begin // @[CSR.scala 50:77]
          mepc <= _GEN_24;
        end
      end
    end
    if (reset) begin // @[CSR.scala 40:23]
      mcause <= 64'h0; // @[CSR.scala 40:23]
    end else if (io_decoderInput_valid) begin // @[CSR.scala 44:31]
      if (!(io_decoderInput_bits_address == 12'hc00 | io_decoderInput_bits_address == 12'hb00)) begin // @[CSR.scala 48:67]
        if (!(io_decoderInput_bits_address == 12'hc02 | io_decoderInput_bits_address == 12'hb02)) begin // @[CSR.scala 50:77]
          mcause <= _GEN_25;
        end
      end
    end
    if (reset) begin // @[CSR.scala 42:24]
      mstatus <= 64'h0; // @[CSR.scala 42:24]
    end else if (io_decoderInput_valid) begin // @[CSR.scala 44:31]
      if (!(io_decoderInput_bits_address == 12'hc00 | io_decoderInput_bits_address == 12'hb00)) begin // @[CSR.scala 48:67]
        if (!(io_decoderInput_bits_address == 12'hc02 | io_decoderInput_bits_address == 12'hb02)) begin // @[CSR.scala 50:77]
          mstatus <= _GEN_26;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  mtvec = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  mepc = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  mcause = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  mstatus = _RAND_3[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CSR_1(
  input         clock,
  input         reset,
  output        io_decoderInput_ready,
  input         io_decoderInput_valid,
  input  [11:0] io_decoderInput_bits_address,
  input  [63:0] io_decoderInput_bits_value,
  input         io_decoderInput_bits_destinationTag_threadId,
  input  [3:0]  io_decoderInput_bits_destinationTag_id,
  input  [1:0]  io_decoderInput_bits_csrAccessType,
  input         io_CSROutput_ready,
  output        io_CSROutput_valid,
  output [63:0] io_CSROutput_bits_value,
  output        io_CSROutput_bits_isError,
  output        io_CSROutput_bits_tag_threadId,
  output [3:0]  io_CSROutput_bits_tag_id,
  output [63:0] io_fetch_mtvec,
  output [63:0] io_fetch_mepc,
  output [63:0] io_fetch_mcause,
  input  [1:0]  io_reorderBuffer_retireCount
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  retireCounter_clock; // @[CSR.scala 32:29]
  wire  retireCounter_reset; // @[CSR.scala 32:29]
  wire [1:0] retireCounter_io_retireInCycle; // @[CSR.scala 32:29]
  wire [63:0] retireCounter_io_count; // @[CSR.scala 32:29]
  wire  cycleCounter_clock; // @[CSR.scala 34:28]
  wire  cycleCounter_reset; // @[CSR.scala 34:28]
  wire [63:0] cycleCounter_count; // @[CSR.scala 34:28]
  reg [63:0] mtvec; // @[CSR.scala 36:22]
  reg [63:0] mepc; // @[CSR.scala 38:21]
  reg [63:0] mcause; // @[CSR.scala 40:23]
  reg [63:0] mstatus; // @[CSR.scala 42:24]
  wire  _T_8 = io_CSROutput_ready & io_CSROutput_valid; // @[CSR.scala 56:31]
  wire [63:0] _mtvec_T_3 = mtvec | io_decoderInput_bits_value; // @[CSR.scala 62:52]
  wire [63:0] _mtvec_T_5 = mtvec & io_decoderInput_bits_value; // @[CSR.scala 63:54]
  wire [63:0] _mtvec_T_7 = 2'h0 == io_decoderInput_bits_csrAccessType ? io_decoderInput_bits_value : 64'h0; // @[Mux.scala 81:58]
  wire [63:0] _mtvec_T_9 = 2'h1 == io_decoderInput_bits_csrAccessType ? _mtvec_T_3 : _mtvec_T_7; // @[Mux.scala 81:58]
  wire [63:0] _mtvec_T_11 = 2'h2 == io_decoderInput_bits_csrAccessType ? _mtvec_T_5 : _mtvec_T_9; // @[Mux.scala 81:58]
  wire [63:0] _GEN_0 = io_CSROutput_ready & io_CSROutput_valid ? _mtvec_T_11 : mtvec; // @[CSR.scala 56:54 57:15 36:22]
  wire [63:0] _mepc_T_3 = mepc | io_decoderInput_bits_value; // @[CSR.scala 75:51]
  wire [63:0] _mepc_T_5 = mepc & io_decoderInput_bits_value; // @[CSR.scala 76:53]
  wire [63:0] _mepc_T_9 = 2'h1 == io_decoderInput_bits_csrAccessType ? _mepc_T_3 : _mtvec_T_7; // @[Mux.scala 81:58]
  wire [63:0] _mepc_T_11 = 2'h2 == io_decoderInput_bits_csrAccessType ? _mepc_T_5 : _mepc_T_9; // @[Mux.scala 81:58]
  wire [63:0] _GEN_1 = _T_8 ? _mepc_T_11 : mepc; // @[CSR.scala 69:54 70:14 38:21]
  wire [63:0] _mcause_T_3 = mcause | io_decoderInput_bits_value; // @[CSR.scala 88:53]
  wire [63:0] _mcause_T_5 = mcause & io_decoderInput_bits_value; // @[CSR.scala 89:55]
  wire [63:0] _mcause_T_9 = 2'h1 == io_decoderInput_bits_csrAccessType ? _mcause_T_3 : _mtvec_T_7; // @[Mux.scala 81:58]
  wire [63:0] _mcause_T_11 = 2'h2 == io_decoderInput_bits_csrAccessType ? _mcause_T_5 : _mcause_T_9; // @[Mux.scala 81:58]
  wire [63:0] _GEN_2 = _T_8 ? _mcause_T_11 : mcause; // @[CSR.scala 82:54 83:16 40:23]
  wire [63:0] _mstatus_T_3 = mstatus | io_decoderInput_bits_value; // @[CSR.scala 101:54]
  wire [63:0] _mstatus_T_5 = mstatus & io_decoderInput_bits_value; // @[CSR.scala 102:56]
  wire [63:0] _mstatus_T_9 = 2'h1 == io_decoderInput_bits_csrAccessType ? _mstatus_T_3 : _mtvec_T_7; // @[Mux.scala 81:58]
  wire [63:0] _mstatus_T_11 = 2'h2 == io_decoderInput_bits_csrAccessType ? _mstatus_T_5 : _mstatus_T_9; // @[Mux.scala 81:58]
  wire [63:0] _GEN_3 = _T_8 ? _mstatus_T_11 : mstatus; // @[CSR.scala 95:54 96:17 42:24]
  wire [63:0] _GEN_4 = io_decoderInput_bits_address == 12'h300 ? mstatus : 64'h0; // @[CSR.scala 26:27 93:45 94:31]
  wire [63:0] _GEN_5 = io_decoderInput_bits_address == 12'h300 ? _GEN_3 : mstatus; // @[CSR.scala 42:24 93:45]
  wire  _GEN_6 = io_decoderInput_bits_address == 12'h300 ? 1'h0 : 1'h1; // @[CSR.scala 27:29 107:33 93:45]
  wire [63:0] _GEN_7 = io_decoderInput_bits_address == 12'h342 ? mcause : _GEN_4; // @[CSR.scala 80:44 81:31]
  wire [63:0] _GEN_8 = io_decoderInput_bits_address == 12'h342 ? _GEN_2 : mcause; // @[CSR.scala 40:23 80:44]
  wire [63:0] _GEN_9 = io_decoderInput_bits_address == 12'h342 ? mstatus : _GEN_5; // @[CSR.scala 42:24 80:44]
  wire  _GEN_10 = io_decoderInput_bits_address == 12'h342 ? 1'h0 : _GEN_6; // @[CSR.scala 27:29 80:44]
  wire [63:0] _GEN_11 = io_decoderInput_bits_address == 12'h341 ? mepc : _GEN_7; // @[CSR.scala 67:42 68:31]
  wire [63:0] _GEN_12 = io_decoderInput_bits_address == 12'h341 ? _GEN_1 : mepc; // @[CSR.scala 38:21 67:42]
  wire [63:0] _GEN_13 = io_decoderInput_bits_address == 12'h341 ? mcause : _GEN_8; // @[CSR.scala 40:23 67:42]
  wire [63:0] _GEN_14 = io_decoderInput_bits_address == 12'h341 ? mstatus : _GEN_9; // @[CSR.scala 42:24 67:42]
  wire  _GEN_15 = io_decoderInput_bits_address == 12'h341 ? 1'h0 : _GEN_10; // @[CSR.scala 27:29 67:42]
  wire [63:0] _GEN_16 = io_decoderInput_bits_address == 12'h305 ? mtvec : _GEN_11; // @[CSR.scala 54:43 55:31]
  wire [63:0] _GEN_17 = io_decoderInput_bits_address == 12'h305 ? _GEN_0 : mtvec; // @[CSR.scala 36:22 54:43]
  wire [63:0] _GEN_18 = io_decoderInput_bits_address == 12'h305 ? mepc : _GEN_12; // @[CSR.scala 38:21 54:43]
  wire [63:0] _GEN_19 = io_decoderInput_bits_address == 12'h305 ? mcause : _GEN_13; // @[CSR.scala 40:23 54:43]
  wire [63:0] _GEN_20 = io_decoderInput_bits_address == 12'h305 ? mstatus : _GEN_14; // @[CSR.scala 42:24 54:43]
  wire  _GEN_21 = io_decoderInput_bits_address == 12'h305 ? 1'h0 : _GEN_15; // @[CSR.scala 27:29 54:43]
  wire [63:0] _GEN_22 = io_decoderInput_bits_address == 12'hf14 ? 64'h1 : _GEN_16; // @[CSR.scala 52:45 53:31]
  wire [63:0] _GEN_23 = io_decoderInput_bits_address == 12'hf14 ? mtvec : _GEN_17; // @[CSR.scala 36:22 52:45]
  wire [63:0] _GEN_24 = io_decoderInput_bits_address == 12'hf14 ? mepc : _GEN_18; // @[CSR.scala 38:21 52:45]
  wire [63:0] _GEN_25 = io_decoderInput_bits_address == 12'hf14 ? mcause : _GEN_19; // @[CSR.scala 40:23 52:45]
  wire [63:0] _GEN_26 = io_decoderInput_bits_address == 12'hf14 ? mstatus : _GEN_20; // @[CSR.scala 42:24 52:45]
  wire  _GEN_27 = io_decoderInput_bits_address == 12'hf14 ? 1'h0 : _GEN_21; // @[CSR.scala 27:29 52:45]
  wire [63:0] _GEN_28 = io_decoderInput_bits_address == 12'hc02 | io_decoderInput_bits_address == 12'hb02 ?
    retireCounter_io_count : _GEN_22; // @[CSR.scala 50:77 51:31]
  wire  _GEN_33 = io_decoderInput_bits_address == 12'hc02 | io_decoderInput_bits_address == 12'hb02 ? 1'h0 : _GEN_27; // @[CSR.scala 27:29 50:77]
  wire [63:0] _GEN_34 = io_decoderInput_bits_address == 12'hc00 | io_decoderInput_bits_address == 12'hb00 ?
    cycleCounter_count : _GEN_28; // @[CSR.scala 48:67 49:31]
  wire  _GEN_39 = io_decoderInput_bits_address == 12'hc00 | io_decoderInput_bits_address == 12'hb00 ? 1'h0 : _GEN_33; // @[CSR.scala 27:29 48:67]
  RetireCounter retireCounter ( // @[CSR.scala 32:29]
    .clock(retireCounter_clock),
    .reset(retireCounter_reset),
    .io_retireInCycle(retireCounter_io_retireInCycle),
    .io_count(retireCounter_io_count)
  );
  CycleCounter cycleCounter ( // @[CSR.scala 34:28]
    .clock(cycleCounter_clock),
    .reset(cycleCounter_reset),
    .count(cycleCounter_count)
  );
  assign io_decoderInput_ready = io_CSROutput_ready; // @[CSR.scala 23:25]
  assign io_CSROutput_valid = io_decoderInput_valid; // @[CSR.scala 24:22 44:31 46:24]
  assign io_CSROutput_bits_value = io_decoderInput_valid ? _GEN_34 : 64'h0; // @[CSR.scala 26:27 44:31]
  assign io_CSROutput_bits_isError = io_decoderInput_valid & _GEN_39; // @[CSR.scala 27:29 44:31]
  assign io_CSROutput_bits_tag_threadId = io_decoderInput_bits_destinationTag_threadId; // @[CSR.scala 25:25]
  assign io_CSROutput_bits_tag_id = io_decoderInput_bits_destinationTag_id; // @[CSR.scala 25:25]
  assign io_fetch_mtvec = mtvec; // @[CSR.scala 37:18]
  assign io_fetch_mepc = mepc; // @[CSR.scala 39:17]
  assign io_fetch_mcause = mcause; // @[CSR.scala 41:19]
  assign retireCounter_clock = clock;
  assign retireCounter_reset = reset;
  assign retireCounter_io_retireInCycle = io_reorderBuffer_retireCount; // @[CSR.scala 33:34]
  assign cycleCounter_clock = clock;
  assign cycleCounter_reset = reset;
  always @(posedge clock) begin
    if (reset) begin // @[CSR.scala 36:22]
      mtvec <= 64'h0; // @[CSR.scala 36:22]
    end else if (io_decoderInput_valid) begin // @[CSR.scala 44:31]
      if (!(io_decoderInput_bits_address == 12'hc00 | io_decoderInput_bits_address == 12'hb00)) begin // @[CSR.scala 48:67]
        if (!(io_decoderInput_bits_address == 12'hc02 | io_decoderInput_bits_address == 12'hb02)) begin // @[CSR.scala 50:77]
          mtvec <= _GEN_23;
        end
      end
    end
    if (reset) begin // @[CSR.scala 38:21]
      mepc <= 64'h0; // @[CSR.scala 38:21]
    end else if (io_decoderInput_valid) begin // @[CSR.scala 44:31]
      if (!(io_decoderInput_bits_address == 12'hc00 | io_decoderInput_bits_address == 12'hb00)) begin // @[CSR.scala 48:67]
        if (!(io_decoderInput_bits_address == 12'hc02 | io_decoderInput_bits_address == 12'hb02)) begin // @[CSR.scala 50:77]
          mepc <= _GEN_24;
        end
      end
    end
    if (reset) begin // @[CSR.scala 40:23]
      mcause <= 64'h0; // @[CSR.scala 40:23]
    end else if (io_decoderInput_valid) begin // @[CSR.scala 44:31]
      if (!(io_decoderInput_bits_address == 12'hc00 | io_decoderInput_bits_address == 12'hb00)) begin // @[CSR.scala 48:67]
        if (!(io_decoderInput_bits_address == 12'hc02 | io_decoderInput_bits_address == 12'hb02)) begin // @[CSR.scala 50:77]
          mcause <= _GEN_25;
        end
      end
    end
    if (reset) begin // @[CSR.scala 42:24]
      mstatus <= 64'h0; // @[CSR.scala 42:24]
    end else if (io_decoderInput_valid) begin // @[CSR.scala 44:31]
      if (!(io_decoderInput_bits_address == 12'hc00 | io_decoderInput_bits_address == 12'hb00)) begin // @[CSR.scala 48:67]
        if (!(io_decoderInput_bits_address == 12'hc02 | io_decoderInput_bits_address == 12'hb02)) begin // @[CSR.scala 50:77]
          mstatus <= _GEN_26;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  mtvec = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  mepc = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  mcause = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  mstatus = _RAND_3[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module B4Processor(
  input         clock,
  input         reset,
  input         axi_writeAddress_ready,
  output        axi_writeAddress_valid,
  output [63:0] axi_writeAddress_bits_ADDR,
  output [7:0]  axi_writeAddress_bits_LEN,
  output [2:0]  axi_writeAddress_bits_SIZE,
  output [1:0]  axi_writeAddress_bits_BURST,
  output        axi_writeAddress_bits_LOCK,
  output [3:0]  axi_writeAddress_bits_CACHE,
  output [2:0]  axi_writeAddress_bits_PROT,
  output [3:0]  axi_writeAddress_bits_QOS,
  output [3:0]  axi_writeAddress_bits_REGION,
  input         axi_write_ready,
  output        axi_write_valid,
  output [63:0] axi_write_bits_DATA,
  output [7:0]  axi_write_bits_STRB,
  output        axi_write_bits_LAST,
  output        axi_writeResponse_ready,
  input         axi_writeResponse_valid,
  input  [1:0]  axi_writeResponse_bits_RESP,
  input         axi_readAddress_ready,
  output        axi_readAddress_valid,
  output [63:0] axi_readAddress_bits_ADDR,
  output [7:0]  axi_readAddress_bits_LEN,
  output [2:0]  axi_readAddress_bits_SIZE,
  output [1:0]  axi_readAddress_bits_BURST,
  output        axi_readAddress_bits_LOCK,
  output [3:0]  axi_readAddress_bits_CACHE,
  output [2:0]  axi_readAddress_bits_PROT,
  output [3:0]  axi_readAddress_bits_QOS,
  output [3:0]  axi_readAddress_bits_REGION,
  output        axi_read_ready,
  input         axi_read_valid,
  input  [63:0] axi_read_bits_DATA,
  input  [1:0]  axi_read_bits_RESP,
  input         axi_read_bits_LAST
);
  wire  instructionCache_0_clock; // @[B4Processor.scala 35:45]
  wire  instructionCache_0_reset; // @[B4Processor.scala 35:45]
  wire  instructionCache_0_io_fetch_0_address_valid; // @[B4Processor.scala 35:45]
  wire [63:0] instructionCache_0_io_fetch_0_address_bits; // @[B4Processor.scala 35:45]
  wire  instructionCache_0_io_fetch_0_output_valid; // @[B4Processor.scala 35:45]
  wire [31:0] instructionCache_0_io_fetch_0_output_bits; // @[B4Processor.scala 35:45]
  wire  instructionCache_0_io_memory_request_ready; // @[B4Processor.scala 35:45]
  wire  instructionCache_0_io_memory_request_valid; // @[B4Processor.scala 35:45]
  wire [63:0] instructionCache_0_io_memory_request_bits_address; // @[B4Processor.scala 35:45]
  wire  instructionCache_0_io_memory_response_valid; // @[B4Processor.scala 35:45]
  wire [63:0] instructionCache_0_io_memory_response_bits_inner; // @[B4Processor.scala 35:45]
  wire  instructionCache_1_clock; // @[B4Processor.scala 35:45]
  wire  instructionCache_1_reset; // @[B4Processor.scala 35:45]
  wire  instructionCache_1_io_fetch_0_address_valid; // @[B4Processor.scala 35:45]
  wire [63:0] instructionCache_1_io_fetch_0_address_bits; // @[B4Processor.scala 35:45]
  wire  instructionCache_1_io_fetch_0_output_valid; // @[B4Processor.scala 35:45]
  wire [31:0] instructionCache_1_io_fetch_0_output_bits; // @[B4Processor.scala 35:45]
  wire  instructionCache_1_io_memory_request_ready; // @[B4Processor.scala 35:45]
  wire  instructionCache_1_io_memory_request_valid; // @[B4Processor.scala 35:45]
  wire [63:0] instructionCache_1_io_memory_request_bits_address; // @[B4Processor.scala 35:45]
  wire  instructionCache_1_io_memory_response_valid; // @[B4Processor.scala 35:45]
  wire [63:0] instructionCache_1_io_memory_response_bits_inner; // @[B4Processor.scala 35:45]
  wire  fetch_0_clock; // @[B4Processor.scala 36:63]
  wire  fetch_0_reset; // @[B4Processor.scala 36:63]
  wire  fetch_0_io_cache_0_address_valid; // @[B4Processor.scala 36:63]
  wire [63:0] fetch_0_io_cache_0_address_bits; // @[B4Processor.scala 36:63]
  wire  fetch_0_io_cache_0_output_valid; // @[B4Processor.scala 36:63]
  wire [31:0] fetch_0_io_cache_0_output_bits; // @[B4Processor.scala 36:63]
  wire  fetch_0_io_reorderBufferEmpty; // @[B4Processor.scala 36:63]
  wire  fetch_0_io_loadStoreQueueEmpty; // @[B4Processor.scala 36:63]
  wire  fetch_0_io_collectedBranchAddresses_addresses_valid; // @[B4Processor.scala 36:63]
  wire  fetch_0_io_collectedBranchAddresses_addresses_bits_threadId; // @[B4Processor.scala 36:63]
  wire [63:0] fetch_0_io_collectedBranchAddresses_addresses_bits_programCounterOffset; // @[B4Processor.scala 36:63]
  wire  fetch_0_io_fetchBuffer_toBuffer_0_ready; // @[B4Processor.scala 36:63]
  wire  fetch_0_io_fetchBuffer_toBuffer_0_valid; // @[B4Processor.scala 36:63]
  wire [31:0] fetch_0_io_fetchBuffer_toBuffer_0_bits_instruction; // @[B4Processor.scala 36:63]
  wire [63:0] fetch_0_io_fetchBuffer_toBuffer_0_bits_programCounter; // @[B4Processor.scala 36:63]
  wire  fetch_0_io_fetchBuffer_empty; // @[B4Processor.scala 36:63]
  wire [63:0] fetch_0_io_csr_mtvec; // @[B4Processor.scala 36:63]
  wire [63:0] fetch_0_io_csr_mepc; // @[B4Processor.scala 36:63]
  wire [63:0] fetch_0_io_csr_mcause; // @[B4Processor.scala 36:63]
  wire  fetch_0_io_csrReservationStationEmpty; // @[B4Processor.scala 36:63]
  wire  fetch_0_io_isError; // @[B4Processor.scala 36:63]
  wire  fetch_1_clock; // @[B4Processor.scala 36:63]
  wire  fetch_1_reset; // @[B4Processor.scala 36:63]
  wire  fetch_1_io_cache_0_address_valid; // @[B4Processor.scala 36:63]
  wire [63:0] fetch_1_io_cache_0_address_bits; // @[B4Processor.scala 36:63]
  wire  fetch_1_io_cache_0_output_valid; // @[B4Processor.scala 36:63]
  wire [31:0] fetch_1_io_cache_0_output_bits; // @[B4Processor.scala 36:63]
  wire  fetch_1_io_reorderBufferEmpty; // @[B4Processor.scala 36:63]
  wire  fetch_1_io_loadStoreQueueEmpty; // @[B4Processor.scala 36:63]
  wire  fetch_1_io_collectedBranchAddresses_addresses_valid; // @[B4Processor.scala 36:63]
  wire  fetch_1_io_collectedBranchAddresses_addresses_bits_threadId; // @[B4Processor.scala 36:63]
  wire [63:0] fetch_1_io_collectedBranchAddresses_addresses_bits_programCounterOffset; // @[B4Processor.scala 36:63]
  wire  fetch_1_io_fetchBuffer_toBuffer_0_ready; // @[B4Processor.scala 36:63]
  wire  fetch_1_io_fetchBuffer_toBuffer_0_valid; // @[B4Processor.scala 36:63]
  wire [31:0] fetch_1_io_fetchBuffer_toBuffer_0_bits_instruction; // @[B4Processor.scala 36:63]
  wire [63:0] fetch_1_io_fetchBuffer_toBuffer_0_bits_programCounter; // @[B4Processor.scala 36:63]
  wire  fetch_1_io_fetchBuffer_empty; // @[B4Processor.scala 36:63]
  wire [63:0] fetch_1_io_csr_mtvec; // @[B4Processor.scala 36:63]
  wire [63:0] fetch_1_io_csr_mepc; // @[B4Processor.scala 36:63]
  wire [63:0] fetch_1_io_csr_mcause; // @[B4Processor.scala 36:63]
  wire  fetch_1_io_csrReservationStationEmpty; // @[B4Processor.scala 36:63]
  wire  fetch_1_io_isError; // @[B4Processor.scala 36:63]
  wire  fetchBuffer_0_clock; // @[B4Processor.scala 38:45]
  wire  fetchBuffer_0_reset; // @[B4Processor.scala 38:45]
  wire  fetchBuffer_0_io_output_0_ready; // @[B4Processor.scala 38:45]
  wire  fetchBuffer_0_io_output_0_valid; // @[B4Processor.scala 38:45]
  wire [31:0] fetchBuffer_0_io_output_0_bits_instruction; // @[B4Processor.scala 38:45]
  wire [63:0] fetchBuffer_0_io_output_0_bits_programCounter; // @[B4Processor.scala 38:45]
  wire  fetchBuffer_0_io_input_toBuffer_0_ready; // @[B4Processor.scala 38:45]
  wire  fetchBuffer_0_io_input_toBuffer_0_valid; // @[B4Processor.scala 38:45]
  wire [31:0] fetchBuffer_0_io_input_toBuffer_0_bits_instruction; // @[B4Processor.scala 38:45]
  wire [63:0] fetchBuffer_0_io_input_toBuffer_0_bits_programCounter; // @[B4Processor.scala 38:45]
  wire  fetchBuffer_0_io_input_empty; // @[B4Processor.scala 38:45]
  wire  fetchBuffer_1_clock; // @[B4Processor.scala 38:45]
  wire  fetchBuffer_1_reset; // @[B4Processor.scala 38:45]
  wire  fetchBuffer_1_io_output_0_ready; // @[B4Processor.scala 38:45]
  wire  fetchBuffer_1_io_output_0_valid; // @[B4Processor.scala 38:45]
  wire [31:0] fetchBuffer_1_io_output_0_bits_instruction; // @[B4Processor.scala 38:45]
  wire [63:0] fetchBuffer_1_io_output_0_bits_programCounter; // @[B4Processor.scala 38:45]
  wire  fetchBuffer_1_io_input_toBuffer_0_ready; // @[B4Processor.scala 38:45]
  wire  fetchBuffer_1_io_input_toBuffer_0_valid; // @[B4Processor.scala 38:45]
  wire [31:0] fetchBuffer_1_io_input_toBuffer_0_bits_instruction; // @[B4Processor.scala 38:45]
  wire [63:0] fetchBuffer_1_io_input_toBuffer_0_bits_programCounter; // @[B4Processor.scala 38:45]
  wire  fetchBuffer_1_io_input_empty; // @[B4Processor.scala 38:45]
  wire  reorderBuffer_0_clock; // @[B4Processor.scala 40:45]
  wire  reorderBuffer_0_reset; // @[B4Processor.scala 40:45]
  wire [4:0] reorderBuffer_0_io_decoders_0_source1_sourceRegister; // @[B4Processor.scala 40:45]
  wire  reorderBuffer_0_io_decoders_0_source1_matchingTag_valid; // @[B4Processor.scala 40:45]
  wire [3:0] reorderBuffer_0_io_decoders_0_source1_matchingTag_bits_id; // @[B4Processor.scala 40:45]
  wire  reorderBuffer_0_io_decoders_0_source1_value_valid; // @[B4Processor.scala 40:45]
  wire [63:0] reorderBuffer_0_io_decoders_0_source1_value_bits; // @[B4Processor.scala 40:45]
  wire [4:0] reorderBuffer_0_io_decoders_0_source2_sourceRegister; // @[B4Processor.scala 40:45]
  wire  reorderBuffer_0_io_decoders_0_source2_matchingTag_valid; // @[B4Processor.scala 40:45]
  wire [3:0] reorderBuffer_0_io_decoders_0_source2_matchingTag_bits_id; // @[B4Processor.scala 40:45]
  wire  reorderBuffer_0_io_decoders_0_source2_value_valid; // @[B4Processor.scala 40:45]
  wire [63:0] reorderBuffer_0_io_decoders_0_source2_value_bits; // @[B4Processor.scala 40:45]
  wire [4:0] reorderBuffer_0_io_decoders_0_destination_destinationRegister; // @[B4Processor.scala 40:45]
  wire [3:0] reorderBuffer_0_io_decoders_0_destination_destinationTag_id; // @[B4Processor.scala 40:45]
  wire  reorderBuffer_0_io_decoders_0_destination_storeSign; // @[B4Processor.scala 40:45]
  wire  reorderBuffer_0_io_decoders_0_ready; // @[B4Processor.scala 40:45]
  wire  reorderBuffer_0_io_decoders_0_valid; // @[B4Processor.scala 40:45]
  wire  reorderBuffer_0_io_collectedOutputs_outputs_valid; // @[B4Processor.scala 40:45]
  wire  reorderBuffer_0_io_collectedOutputs_outputs_bits_resultType; // @[B4Processor.scala 40:45]
  wire [63:0] reorderBuffer_0_io_collectedOutputs_outputs_bits_value; // @[B4Processor.scala 40:45]
  wire  reorderBuffer_0_io_collectedOutputs_outputs_bits_isError; // @[B4Processor.scala 40:45]
  wire  reorderBuffer_0_io_collectedOutputs_outputs_bits_tag_threadId; // @[B4Processor.scala 40:45]
  wire [3:0] reorderBuffer_0_io_collectedOutputs_outputs_bits_tag_id; // @[B4Processor.scala 40:45]
  wire  reorderBuffer_0_io_registerFile_0_valid; // @[B4Processor.scala 40:45]
  wire [4:0] reorderBuffer_0_io_registerFile_0_bits_destinationRegister; // @[B4Processor.scala 40:45]
  wire [63:0] reorderBuffer_0_io_registerFile_0_bits_value; // @[B4Processor.scala 40:45]
  wire  reorderBuffer_0_io_registerFile_1_valid; // @[B4Processor.scala 40:45]
  wire [4:0] reorderBuffer_0_io_registerFile_1_bits_destinationRegister; // @[B4Processor.scala 40:45]
  wire [63:0] reorderBuffer_0_io_registerFile_1_bits_value; // @[B4Processor.scala 40:45]
  wire  reorderBuffer_0_io_registerFile_2_valid; // @[B4Processor.scala 40:45]
  wire [4:0] reorderBuffer_0_io_registerFile_2_bits_destinationRegister; // @[B4Processor.scala 40:45]
  wire [63:0] reorderBuffer_0_io_registerFile_2_bits_value; // @[B4Processor.scala 40:45]
  wire  reorderBuffer_0_io_registerFile_3_valid; // @[B4Processor.scala 40:45]
  wire [4:0] reorderBuffer_0_io_registerFile_3_bits_destinationRegister; // @[B4Processor.scala 40:45]
  wire [63:0] reorderBuffer_0_io_registerFile_3_bits_value; // @[B4Processor.scala 40:45]
  wire  reorderBuffer_0_io_loadStoreQueue_0_valid; // @[B4Processor.scala 40:45]
  wire [3:0] reorderBuffer_0_io_loadStoreQueue_0_bits_destinationTag_id; // @[B4Processor.scala 40:45]
  wire  reorderBuffer_0_io_loadStoreQueue_1_valid; // @[B4Processor.scala 40:45]
  wire [3:0] reorderBuffer_0_io_loadStoreQueue_1_bits_destinationTag_id; // @[B4Processor.scala 40:45]
  wire  reorderBuffer_0_io_loadStoreQueue_2_valid; // @[B4Processor.scala 40:45]
  wire [3:0] reorderBuffer_0_io_loadStoreQueue_2_bits_destinationTag_id; // @[B4Processor.scala 40:45]
  wire  reorderBuffer_0_io_loadStoreQueue_3_valid; // @[B4Processor.scala 40:45]
  wire [3:0] reorderBuffer_0_io_loadStoreQueue_3_bits_destinationTag_id; // @[B4Processor.scala 40:45]
  wire  reorderBuffer_0_io_isEmpty; // @[B4Processor.scala 40:45]
  wire [1:0] reorderBuffer_0_io_csr_retireCount; // @[B4Processor.scala 40:45]
  wire  reorderBuffer_0_io_isError; // @[B4Processor.scala 40:45]
  wire  reorderBuffer_1_clock; // @[B4Processor.scala 40:45]
  wire  reorderBuffer_1_reset; // @[B4Processor.scala 40:45]
  wire [4:0] reorderBuffer_1_io_decoders_0_source1_sourceRegister; // @[B4Processor.scala 40:45]
  wire  reorderBuffer_1_io_decoders_0_source1_matchingTag_valid; // @[B4Processor.scala 40:45]
  wire [3:0] reorderBuffer_1_io_decoders_0_source1_matchingTag_bits_id; // @[B4Processor.scala 40:45]
  wire  reorderBuffer_1_io_decoders_0_source1_value_valid; // @[B4Processor.scala 40:45]
  wire [63:0] reorderBuffer_1_io_decoders_0_source1_value_bits; // @[B4Processor.scala 40:45]
  wire [4:0] reorderBuffer_1_io_decoders_0_source2_sourceRegister; // @[B4Processor.scala 40:45]
  wire  reorderBuffer_1_io_decoders_0_source2_matchingTag_valid; // @[B4Processor.scala 40:45]
  wire [3:0] reorderBuffer_1_io_decoders_0_source2_matchingTag_bits_id; // @[B4Processor.scala 40:45]
  wire  reorderBuffer_1_io_decoders_0_source2_value_valid; // @[B4Processor.scala 40:45]
  wire [63:0] reorderBuffer_1_io_decoders_0_source2_value_bits; // @[B4Processor.scala 40:45]
  wire [4:0] reorderBuffer_1_io_decoders_0_destination_destinationRegister; // @[B4Processor.scala 40:45]
  wire [3:0] reorderBuffer_1_io_decoders_0_destination_destinationTag_id; // @[B4Processor.scala 40:45]
  wire  reorderBuffer_1_io_decoders_0_destination_storeSign; // @[B4Processor.scala 40:45]
  wire  reorderBuffer_1_io_decoders_0_ready; // @[B4Processor.scala 40:45]
  wire  reorderBuffer_1_io_decoders_0_valid; // @[B4Processor.scala 40:45]
  wire  reorderBuffer_1_io_collectedOutputs_outputs_valid; // @[B4Processor.scala 40:45]
  wire  reorderBuffer_1_io_collectedOutputs_outputs_bits_resultType; // @[B4Processor.scala 40:45]
  wire [63:0] reorderBuffer_1_io_collectedOutputs_outputs_bits_value; // @[B4Processor.scala 40:45]
  wire  reorderBuffer_1_io_collectedOutputs_outputs_bits_isError; // @[B4Processor.scala 40:45]
  wire  reorderBuffer_1_io_collectedOutputs_outputs_bits_tag_threadId; // @[B4Processor.scala 40:45]
  wire [3:0] reorderBuffer_1_io_collectedOutputs_outputs_bits_tag_id; // @[B4Processor.scala 40:45]
  wire  reorderBuffer_1_io_registerFile_0_valid; // @[B4Processor.scala 40:45]
  wire [4:0] reorderBuffer_1_io_registerFile_0_bits_destinationRegister; // @[B4Processor.scala 40:45]
  wire [63:0] reorderBuffer_1_io_registerFile_0_bits_value; // @[B4Processor.scala 40:45]
  wire  reorderBuffer_1_io_registerFile_1_valid; // @[B4Processor.scala 40:45]
  wire [4:0] reorderBuffer_1_io_registerFile_1_bits_destinationRegister; // @[B4Processor.scala 40:45]
  wire [63:0] reorderBuffer_1_io_registerFile_1_bits_value; // @[B4Processor.scala 40:45]
  wire  reorderBuffer_1_io_registerFile_2_valid; // @[B4Processor.scala 40:45]
  wire [4:0] reorderBuffer_1_io_registerFile_2_bits_destinationRegister; // @[B4Processor.scala 40:45]
  wire [63:0] reorderBuffer_1_io_registerFile_2_bits_value; // @[B4Processor.scala 40:45]
  wire  reorderBuffer_1_io_registerFile_3_valid; // @[B4Processor.scala 40:45]
  wire [4:0] reorderBuffer_1_io_registerFile_3_bits_destinationRegister; // @[B4Processor.scala 40:45]
  wire [63:0] reorderBuffer_1_io_registerFile_3_bits_value; // @[B4Processor.scala 40:45]
  wire  reorderBuffer_1_io_loadStoreQueue_0_valid; // @[B4Processor.scala 40:45]
  wire [3:0] reorderBuffer_1_io_loadStoreQueue_0_bits_destinationTag_id; // @[B4Processor.scala 40:45]
  wire  reorderBuffer_1_io_loadStoreQueue_1_valid; // @[B4Processor.scala 40:45]
  wire [3:0] reorderBuffer_1_io_loadStoreQueue_1_bits_destinationTag_id; // @[B4Processor.scala 40:45]
  wire  reorderBuffer_1_io_loadStoreQueue_2_valid; // @[B4Processor.scala 40:45]
  wire [3:0] reorderBuffer_1_io_loadStoreQueue_2_bits_destinationTag_id; // @[B4Processor.scala 40:45]
  wire  reorderBuffer_1_io_loadStoreQueue_3_valid; // @[B4Processor.scala 40:45]
  wire [3:0] reorderBuffer_1_io_loadStoreQueue_3_bits_destinationTag_id; // @[B4Processor.scala 40:45]
  wire  reorderBuffer_1_io_isEmpty; // @[B4Processor.scala 40:45]
  wire [1:0] reorderBuffer_1_io_csr_retireCount; // @[B4Processor.scala 40:45]
  wire  reorderBuffer_1_io_isError; // @[B4Processor.scala 40:45]
  wire  registerFile_0_clock; // @[B4Processor.scala 42:45]
  wire  registerFile_0_reset; // @[B4Processor.scala 42:45]
  wire [4:0] registerFile_0_io_decoders_0_sourceRegister1; // @[B4Processor.scala 42:45]
  wire [4:0] registerFile_0_io_decoders_0_sourceRegister2; // @[B4Processor.scala 42:45]
  wire [63:0] registerFile_0_io_decoders_0_value1; // @[B4Processor.scala 42:45]
  wire [63:0] registerFile_0_io_decoders_0_value2; // @[B4Processor.scala 42:45]
  wire  registerFile_0_io_reorderBuffer_0_valid; // @[B4Processor.scala 42:45]
  wire [4:0] registerFile_0_io_reorderBuffer_0_bits_destinationRegister; // @[B4Processor.scala 42:45]
  wire [63:0] registerFile_0_io_reorderBuffer_0_bits_value; // @[B4Processor.scala 42:45]
  wire  registerFile_0_io_reorderBuffer_1_valid; // @[B4Processor.scala 42:45]
  wire [4:0] registerFile_0_io_reorderBuffer_1_bits_destinationRegister; // @[B4Processor.scala 42:45]
  wire [63:0] registerFile_0_io_reorderBuffer_1_bits_value; // @[B4Processor.scala 42:45]
  wire  registerFile_0_io_reorderBuffer_2_valid; // @[B4Processor.scala 42:45]
  wire [4:0] registerFile_0_io_reorderBuffer_2_bits_destinationRegister; // @[B4Processor.scala 42:45]
  wire [63:0] registerFile_0_io_reorderBuffer_2_bits_value; // @[B4Processor.scala 42:45]
  wire  registerFile_0_io_reorderBuffer_3_valid; // @[B4Processor.scala 42:45]
  wire [4:0] registerFile_0_io_reorderBuffer_3_bits_destinationRegister; // @[B4Processor.scala 42:45]
  wire [63:0] registerFile_0_io_reorderBuffer_3_bits_value; // @[B4Processor.scala 42:45]
  wire  registerFile_1_clock; // @[B4Processor.scala 42:45]
  wire  registerFile_1_reset; // @[B4Processor.scala 42:45]
  wire [4:0] registerFile_1_io_decoders_0_sourceRegister1; // @[B4Processor.scala 42:45]
  wire [4:0] registerFile_1_io_decoders_0_sourceRegister2; // @[B4Processor.scala 42:45]
  wire [63:0] registerFile_1_io_decoders_0_value1; // @[B4Processor.scala 42:45]
  wire [63:0] registerFile_1_io_decoders_0_value2; // @[B4Processor.scala 42:45]
  wire  registerFile_1_io_reorderBuffer_0_valid; // @[B4Processor.scala 42:45]
  wire [4:0] registerFile_1_io_reorderBuffer_0_bits_destinationRegister; // @[B4Processor.scala 42:45]
  wire [63:0] registerFile_1_io_reorderBuffer_0_bits_value; // @[B4Processor.scala 42:45]
  wire  registerFile_1_io_reorderBuffer_1_valid; // @[B4Processor.scala 42:45]
  wire [4:0] registerFile_1_io_reorderBuffer_1_bits_destinationRegister; // @[B4Processor.scala 42:45]
  wire [63:0] registerFile_1_io_reorderBuffer_1_bits_value; // @[B4Processor.scala 42:45]
  wire  registerFile_1_io_reorderBuffer_2_valid; // @[B4Processor.scala 42:45]
  wire [4:0] registerFile_1_io_reorderBuffer_2_bits_destinationRegister; // @[B4Processor.scala 42:45]
  wire [63:0] registerFile_1_io_reorderBuffer_2_bits_value; // @[B4Processor.scala 42:45]
  wire  registerFile_1_io_reorderBuffer_3_valid; // @[B4Processor.scala 42:45]
  wire [4:0] registerFile_1_io_reorderBuffer_3_bits_destinationRegister; // @[B4Processor.scala 42:45]
  wire [63:0] registerFile_1_io_reorderBuffer_3_bits_value; // @[B4Processor.scala 42:45]
  wire  loadStoreQueue_0_clock; // @[B4Processor.scala 44:45]
  wire  loadStoreQueue_0_reset; // @[B4Processor.scala 44:45]
  wire  loadStoreQueue_0_io_decoders_0_ready; // @[B4Processor.scala 44:45]
  wire  loadStoreQueue_0_io_decoders_0_valid; // @[B4Processor.scala 44:45]
  wire  loadStoreQueue_0_io_decoders_0_bits_accessInfo_accessType; // @[B4Processor.scala 44:45]
  wire  loadStoreQueue_0_io_decoders_0_bits_accessInfo_signed; // @[B4Processor.scala 44:45]
  wire [1:0] loadStoreQueue_0_io_decoders_0_bits_accessInfo_accessWidth; // @[B4Processor.scala 44:45]
  wire  loadStoreQueue_0_io_decoders_0_bits_addressAndLoadResultTag_threadId; // @[B4Processor.scala 44:45]
  wire [3:0] loadStoreQueue_0_io_decoders_0_bits_addressAndLoadResultTag_id; // @[B4Processor.scala 44:45]
  wire [63:0] loadStoreQueue_0_io_decoders_0_bits_address; // @[B4Processor.scala 44:45]
  wire  loadStoreQueue_0_io_decoders_0_bits_addressValid; // @[B4Processor.scala 44:45]
  wire  loadStoreQueue_0_io_decoders_0_bits_storeDataTag_threadId; // @[B4Processor.scala 44:45]
  wire [3:0] loadStoreQueue_0_io_decoders_0_bits_storeDataTag_id; // @[B4Processor.scala 44:45]
  wire [63:0] loadStoreQueue_0_io_decoders_0_bits_storeData; // @[B4Processor.scala 44:45]
  wire  loadStoreQueue_0_io_decoders_0_bits_storeDataValid; // @[B4Processor.scala 44:45]
  wire  loadStoreQueue_0_io_outputCollector_outputs_valid; // @[B4Processor.scala 44:45]
  wire  loadStoreQueue_0_io_outputCollector_outputs_bits_resultType; // @[B4Processor.scala 44:45]
  wire [63:0] loadStoreQueue_0_io_outputCollector_outputs_bits_value; // @[B4Processor.scala 44:45]
  wire  loadStoreQueue_0_io_outputCollector_outputs_bits_tag_threadId; // @[B4Processor.scala 44:45]
  wire [3:0] loadStoreQueue_0_io_outputCollector_outputs_bits_tag_id; // @[B4Processor.scala 44:45]
  wire  loadStoreQueue_0_io_reorderBuffer_0_valid; // @[B4Processor.scala 44:45]
  wire  loadStoreQueue_0_io_reorderBuffer_0_bits_destinationTag_threadId; // @[B4Processor.scala 44:45]
  wire [3:0] loadStoreQueue_0_io_reorderBuffer_0_bits_destinationTag_id; // @[B4Processor.scala 44:45]
  wire  loadStoreQueue_0_io_reorderBuffer_1_valid; // @[B4Processor.scala 44:45]
  wire  loadStoreQueue_0_io_reorderBuffer_1_bits_destinationTag_threadId; // @[B4Processor.scala 44:45]
  wire [3:0] loadStoreQueue_0_io_reorderBuffer_1_bits_destinationTag_id; // @[B4Processor.scala 44:45]
  wire  loadStoreQueue_0_io_reorderBuffer_2_valid; // @[B4Processor.scala 44:45]
  wire  loadStoreQueue_0_io_reorderBuffer_2_bits_destinationTag_threadId; // @[B4Processor.scala 44:45]
  wire [3:0] loadStoreQueue_0_io_reorderBuffer_2_bits_destinationTag_id; // @[B4Processor.scala 44:45]
  wire  loadStoreQueue_0_io_reorderBuffer_3_valid; // @[B4Processor.scala 44:45]
  wire  loadStoreQueue_0_io_reorderBuffer_3_bits_destinationTag_threadId; // @[B4Processor.scala 44:45]
  wire [3:0] loadStoreQueue_0_io_reorderBuffer_3_bits_destinationTag_id; // @[B4Processor.scala 44:45]
  wire  loadStoreQueue_0_io_memory_ready; // @[B4Processor.scala 44:45]
  wire  loadStoreQueue_0_io_memory_valid; // @[B4Processor.scala 44:45]
  wire [63:0] loadStoreQueue_0_io_memory_bits_address; // @[B4Processor.scala 44:45]
  wire  loadStoreQueue_0_io_memory_bits_tag_threadId; // @[B4Processor.scala 44:45]
  wire [3:0] loadStoreQueue_0_io_memory_bits_tag_id; // @[B4Processor.scala 44:45]
  wire [63:0] loadStoreQueue_0_io_memory_bits_data; // @[B4Processor.scala 44:45]
  wire  loadStoreQueue_0_io_memory_bits_accessInfo_accessType; // @[B4Processor.scala 44:45]
  wire  loadStoreQueue_0_io_memory_bits_accessInfo_signed; // @[B4Processor.scala 44:45]
  wire [1:0] loadStoreQueue_0_io_memory_bits_accessInfo_accessWidth; // @[B4Processor.scala 44:45]
  wire  loadStoreQueue_0_io_isEmpty; // @[B4Processor.scala 44:45]
  wire  loadStoreQueue_1_clock; // @[B4Processor.scala 44:45]
  wire  loadStoreQueue_1_reset; // @[B4Processor.scala 44:45]
  wire  loadStoreQueue_1_io_decoders_0_ready; // @[B4Processor.scala 44:45]
  wire  loadStoreQueue_1_io_decoders_0_valid; // @[B4Processor.scala 44:45]
  wire  loadStoreQueue_1_io_decoders_0_bits_accessInfo_accessType; // @[B4Processor.scala 44:45]
  wire  loadStoreQueue_1_io_decoders_0_bits_accessInfo_signed; // @[B4Processor.scala 44:45]
  wire [1:0] loadStoreQueue_1_io_decoders_0_bits_accessInfo_accessWidth; // @[B4Processor.scala 44:45]
  wire  loadStoreQueue_1_io_decoders_0_bits_addressAndLoadResultTag_threadId; // @[B4Processor.scala 44:45]
  wire [3:0] loadStoreQueue_1_io_decoders_0_bits_addressAndLoadResultTag_id; // @[B4Processor.scala 44:45]
  wire [63:0] loadStoreQueue_1_io_decoders_0_bits_address; // @[B4Processor.scala 44:45]
  wire  loadStoreQueue_1_io_decoders_0_bits_addressValid; // @[B4Processor.scala 44:45]
  wire  loadStoreQueue_1_io_decoders_0_bits_storeDataTag_threadId; // @[B4Processor.scala 44:45]
  wire [3:0] loadStoreQueue_1_io_decoders_0_bits_storeDataTag_id; // @[B4Processor.scala 44:45]
  wire [63:0] loadStoreQueue_1_io_decoders_0_bits_storeData; // @[B4Processor.scala 44:45]
  wire  loadStoreQueue_1_io_decoders_0_bits_storeDataValid; // @[B4Processor.scala 44:45]
  wire  loadStoreQueue_1_io_outputCollector_outputs_valid; // @[B4Processor.scala 44:45]
  wire  loadStoreQueue_1_io_outputCollector_outputs_bits_resultType; // @[B4Processor.scala 44:45]
  wire [63:0] loadStoreQueue_1_io_outputCollector_outputs_bits_value; // @[B4Processor.scala 44:45]
  wire  loadStoreQueue_1_io_outputCollector_outputs_bits_tag_threadId; // @[B4Processor.scala 44:45]
  wire [3:0] loadStoreQueue_1_io_outputCollector_outputs_bits_tag_id; // @[B4Processor.scala 44:45]
  wire  loadStoreQueue_1_io_reorderBuffer_0_valid; // @[B4Processor.scala 44:45]
  wire  loadStoreQueue_1_io_reorderBuffer_0_bits_destinationTag_threadId; // @[B4Processor.scala 44:45]
  wire [3:0] loadStoreQueue_1_io_reorderBuffer_0_bits_destinationTag_id; // @[B4Processor.scala 44:45]
  wire  loadStoreQueue_1_io_reorderBuffer_1_valid; // @[B4Processor.scala 44:45]
  wire  loadStoreQueue_1_io_reorderBuffer_1_bits_destinationTag_threadId; // @[B4Processor.scala 44:45]
  wire [3:0] loadStoreQueue_1_io_reorderBuffer_1_bits_destinationTag_id; // @[B4Processor.scala 44:45]
  wire  loadStoreQueue_1_io_reorderBuffer_2_valid; // @[B4Processor.scala 44:45]
  wire  loadStoreQueue_1_io_reorderBuffer_2_bits_destinationTag_threadId; // @[B4Processor.scala 44:45]
  wire [3:0] loadStoreQueue_1_io_reorderBuffer_2_bits_destinationTag_id; // @[B4Processor.scala 44:45]
  wire  loadStoreQueue_1_io_reorderBuffer_3_valid; // @[B4Processor.scala 44:45]
  wire  loadStoreQueue_1_io_reorderBuffer_3_bits_destinationTag_threadId; // @[B4Processor.scala 44:45]
  wire [3:0] loadStoreQueue_1_io_reorderBuffer_3_bits_destinationTag_id; // @[B4Processor.scala 44:45]
  wire  loadStoreQueue_1_io_memory_ready; // @[B4Processor.scala 44:45]
  wire  loadStoreQueue_1_io_memory_valid; // @[B4Processor.scala 44:45]
  wire [63:0] loadStoreQueue_1_io_memory_bits_address; // @[B4Processor.scala 44:45]
  wire  loadStoreQueue_1_io_memory_bits_tag_threadId; // @[B4Processor.scala 44:45]
  wire [3:0] loadStoreQueue_1_io_memory_bits_tag_id; // @[B4Processor.scala 44:45]
  wire [63:0] loadStoreQueue_1_io_memory_bits_data; // @[B4Processor.scala 44:45]
  wire  loadStoreQueue_1_io_memory_bits_accessInfo_accessType; // @[B4Processor.scala 44:45]
  wire  loadStoreQueue_1_io_memory_bits_accessInfo_signed; // @[B4Processor.scala 44:45]
  wire [1:0] loadStoreQueue_1_io_memory_bits_accessInfo_accessWidth; // @[B4Processor.scala 44:45]
  wire  loadStoreQueue_1_io_isEmpty; // @[B4Processor.scala 44:45]
  wire  dataMemoryBuffer_clock; // @[B4Processor.scala 45:40]
  wire  dataMemoryBuffer_reset; // @[B4Processor.scala 45:40]
  wire  dataMemoryBuffer_io_dataIn_0_ready; // @[B4Processor.scala 45:40]
  wire  dataMemoryBuffer_io_dataIn_0_valid; // @[B4Processor.scala 45:40]
  wire [63:0] dataMemoryBuffer_io_dataIn_0_bits_address; // @[B4Processor.scala 45:40]
  wire  dataMemoryBuffer_io_dataIn_0_bits_tag_threadId; // @[B4Processor.scala 45:40]
  wire [3:0] dataMemoryBuffer_io_dataIn_0_bits_tag_id; // @[B4Processor.scala 45:40]
  wire [63:0] dataMemoryBuffer_io_dataIn_0_bits_data; // @[B4Processor.scala 45:40]
  wire  dataMemoryBuffer_io_dataIn_0_bits_accessInfo_accessType; // @[B4Processor.scala 45:40]
  wire  dataMemoryBuffer_io_dataIn_0_bits_accessInfo_signed; // @[B4Processor.scala 45:40]
  wire [1:0] dataMemoryBuffer_io_dataIn_0_bits_accessInfo_accessWidth; // @[B4Processor.scala 45:40]
  wire  dataMemoryBuffer_io_dataIn_1_ready; // @[B4Processor.scala 45:40]
  wire  dataMemoryBuffer_io_dataIn_1_valid; // @[B4Processor.scala 45:40]
  wire [63:0] dataMemoryBuffer_io_dataIn_1_bits_address; // @[B4Processor.scala 45:40]
  wire  dataMemoryBuffer_io_dataIn_1_bits_tag_threadId; // @[B4Processor.scala 45:40]
  wire [3:0] dataMemoryBuffer_io_dataIn_1_bits_tag_id; // @[B4Processor.scala 45:40]
  wire [63:0] dataMemoryBuffer_io_dataIn_1_bits_data; // @[B4Processor.scala 45:40]
  wire  dataMemoryBuffer_io_dataIn_1_bits_accessInfo_accessType; // @[B4Processor.scala 45:40]
  wire  dataMemoryBuffer_io_dataIn_1_bits_accessInfo_signed; // @[B4Processor.scala 45:40]
  wire [1:0] dataMemoryBuffer_io_dataIn_1_bits_accessInfo_accessWidth; // @[B4Processor.scala 45:40]
  wire  dataMemoryBuffer_io_dataReadRequest_ready; // @[B4Processor.scala 45:40]
  wire  dataMemoryBuffer_io_dataReadRequest_valid; // @[B4Processor.scala 45:40]
  wire [63:0] dataMemoryBuffer_io_dataReadRequest_bits_address; // @[B4Processor.scala 45:40]
  wire [1:0] dataMemoryBuffer_io_dataReadRequest_bits_size; // @[B4Processor.scala 45:40]
  wire  dataMemoryBuffer_io_dataReadRequest_bits_signed; // @[B4Processor.scala 45:40]
  wire  dataMemoryBuffer_io_dataReadRequest_bits_outputTag_threadId; // @[B4Processor.scala 45:40]
  wire [3:0] dataMemoryBuffer_io_dataReadRequest_bits_outputTag_id; // @[B4Processor.scala 45:40]
  wire  dataMemoryBuffer_io_dataWriteRequest_ready; // @[B4Processor.scala 45:40]
  wire  dataMemoryBuffer_io_dataWriteRequest_valid; // @[B4Processor.scala 45:40]
  wire [63:0] dataMemoryBuffer_io_dataWriteRequest_bits_address; // @[B4Processor.scala 45:40]
  wire [63:0] dataMemoryBuffer_io_dataWriteRequest_bits_data; // @[B4Processor.scala 45:40]
  wire [7:0] dataMemoryBuffer_io_dataWriteRequest_bits_mask; // @[B4Processor.scala 45:40]
  wire  outputCollector_clock; // @[B4Processor.scala 47:31]
  wire  outputCollector_reset; // @[B4Processor.scala 47:31]
  wire  outputCollector_io_outputs_0_outputs_valid; // @[B4Processor.scala 47:31]
  wire  outputCollector_io_outputs_0_outputs_bits_resultType; // @[B4Processor.scala 47:31]
  wire [63:0] outputCollector_io_outputs_0_outputs_bits_value; // @[B4Processor.scala 47:31]
  wire  outputCollector_io_outputs_0_outputs_bits_isError; // @[B4Processor.scala 47:31]
  wire  outputCollector_io_outputs_0_outputs_bits_tag_threadId; // @[B4Processor.scala 47:31]
  wire [3:0] outputCollector_io_outputs_0_outputs_bits_tag_id; // @[B4Processor.scala 47:31]
  wire  outputCollector_io_outputs_1_outputs_valid; // @[B4Processor.scala 47:31]
  wire  outputCollector_io_outputs_1_outputs_bits_resultType; // @[B4Processor.scala 47:31]
  wire [63:0] outputCollector_io_outputs_1_outputs_bits_value; // @[B4Processor.scala 47:31]
  wire  outputCollector_io_outputs_1_outputs_bits_isError; // @[B4Processor.scala 47:31]
  wire  outputCollector_io_outputs_1_outputs_bits_tag_threadId; // @[B4Processor.scala 47:31]
  wire [3:0] outputCollector_io_outputs_1_outputs_bits_tag_id; // @[B4Processor.scala 47:31]
  wire  outputCollector_io_executor_0_ready; // @[B4Processor.scala 47:31]
  wire  outputCollector_io_executor_0_valid; // @[B4Processor.scala 47:31]
  wire  outputCollector_io_executor_0_bits_resultType; // @[B4Processor.scala 47:31]
  wire [63:0] outputCollector_io_executor_0_bits_value; // @[B4Processor.scala 47:31]
  wire  outputCollector_io_executor_0_bits_tag_threadId; // @[B4Processor.scala 47:31]
  wire [3:0] outputCollector_io_executor_0_bits_tag_id; // @[B4Processor.scala 47:31]
  wire  outputCollector_io_executor_1_ready; // @[B4Processor.scala 47:31]
  wire  outputCollector_io_executor_1_valid; // @[B4Processor.scala 47:31]
  wire  outputCollector_io_executor_1_bits_resultType; // @[B4Processor.scala 47:31]
  wire [63:0] outputCollector_io_executor_1_bits_value; // @[B4Processor.scala 47:31]
  wire  outputCollector_io_executor_1_bits_tag_threadId; // @[B4Processor.scala 47:31]
  wire [3:0] outputCollector_io_executor_1_bits_tag_id; // @[B4Processor.scala 47:31]
  wire  outputCollector_io_dataMemory_ready; // @[B4Processor.scala 47:31]
  wire  outputCollector_io_dataMemory_valid; // @[B4Processor.scala 47:31]
  wire [63:0] outputCollector_io_dataMemory_bits_value; // @[B4Processor.scala 47:31]
  wire  outputCollector_io_dataMemory_bits_isError; // @[B4Processor.scala 47:31]
  wire  outputCollector_io_dataMemory_bits_tag_threadId; // @[B4Processor.scala 47:31]
  wire [3:0] outputCollector_io_dataMemory_bits_tag_id; // @[B4Processor.scala 47:31]
  wire  outputCollector_io_csr_0_ready; // @[B4Processor.scala 47:31]
  wire  outputCollector_io_csr_0_valid; // @[B4Processor.scala 47:31]
  wire [63:0] outputCollector_io_csr_0_bits_value; // @[B4Processor.scala 47:31]
  wire  outputCollector_io_csr_0_bits_isError; // @[B4Processor.scala 47:31]
  wire  outputCollector_io_csr_0_bits_tag_threadId; // @[B4Processor.scala 47:31]
  wire [3:0] outputCollector_io_csr_0_bits_tag_id; // @[B4Processor.scala 47:31]
  wire  outputCollector_io_csr_1_ready; // @[B4Processor.scala 47:31]
  wire  outputCollector_io_csr_1_valid; // @[B4Processor.scala 47:31]
  wire [63:0] outputCollector_io_csr_1_bits_value; // @[B4Processor.scala 47:31]
  wire  outputCollector_io_csr_1_bits_isError; // @[B4Processor.scala 47:31]
  wire  outputCollector_io_csr_1_bits_tag_threadId; // @[B4Processor.scala 47:31]
  wire [3:0] outputCollector_io_csr_1_bits_tag_id; // @[B4Processor.scala 47:31]
  wire  outputCollector_io_isError_0; // @[B4Processor.scala 47:31]
  wire  outputCollector_io_isError_1; // @[B4Processor.scala 47:31]
  wire  branchAddressCollector_clock; // @[B4Processor.scala 48:46]
  wire  branchAddressCollector_reset; // @[B4Processor.scala 48:46]
  wire  branchAddressCollector_io_fetch_0_addresses_valid; // @[B4Processor.scala 48:46]
  wire  branchAddressCollector_io_fetch_0_addresses_bits_threadId; // @[B4Processor.scala 48:46]
  wire [63:0] branchAddressCollector_io_fetch_0_addresses_bits_programCounterOffset; // @[B4Processor.scala 48:46]
  wire  branchAddressCollector_io_fetch_1_addresses_valid; // @[B4Processor.scala 48:46]
  wire  branchAddressCollector_io_fetch_1_addresses_bits_threadId; // @[B4Processor.scala 48:46]
  wire [63:0] branchAddressCollector_io_fetch_1_addresses_bits_programCounterOffset; // @[B4Processor.scala 48:46]
  wire  branchAddressCollector_io_executor_0_ready; // @[B4Processor.scala 48:46]
  wire  branchAddressCollector_io_executor_0_valid; // @[B4Processor.scala 48:46]
  wire  branchAddressCollector_io_executor_0_bits_threadId; // @[B4Processor.scala 48:46]
  wire [63:0] branchAddressCollector_io_executor_0_bits_programCounterOffset; // @[B4Processor.scala 48:46]
  wire  branchAddressCollector_io_executor_1_ready; // @[B4Processor.scala 48:46]
  wire  branchAddressCollector_io_executor_1_valid; // @[B4Processor.scala 48:46]
  wire  branchAddressCollector_io_executor_1_bits_threadId; // @[B4Processor.scala 48:46]
  wire [63:0] branchAddressCollector_io_executor_1_bits_programCounterOffset; // @[B4Processor.scala 48:46]
  wire  branchAddressCollector_io_isError_0; // @[B4Processor.scala 48:46]
  wire  branchAddressCollector_io_isError_1; // @[B4Processor.scala 48:46]
  wire  uncompresser_0_0_io_fetch_ready; // @[B4Processor.scala 51:45]
  wire  uncompresser_0_0_io_fetch_valid; // @[B4Processor.scala 51:45]
  wire [31:0] uncompresser_0_0_io_fetch_bits_instruction; // @[B4Processor.scala 51:45]
  wire [63:0] uncompresser_0_0_io_fetch_bits_programCounter; // @[B4Processor.scala 51:45]
  wire  uncompresser_0_0_io_decoder_ready; // @[B4Processor.scala 51:45]
  wire  uncompresser_0_0_io_decoder_valid; // @[B4Processor.scala 51:45]
  wire [31:0] uncompresser_0_0_io_decoder_bits_instruction; // @[B4Processor.scala 51:45]
  wire [63:0] uncompresser_0_0_io_decoder_bits_programCounter; // @[B4Processor.scala 51:45]
  wire  uncompresser_0_0_io_decoder_bits_wasCompressed; // @[B4Processor.scala 51:45]
  wire  uncompresser_1_0_io_fetch_ready; // @[B4Processor.scala 51:45]
  wire  uncompresser_1_0_io_fetch_valid; // @[B4Processor.scala 51:45]
  wire [31:0] uncompresser_1_0_io_fetch_bits_instruction; // @[B4Processor.scala 51:45]
  wire [63:0] uncompresser_1_0_io_fetch_bits_programCounter; // @[B4Processor.scala 51:45]
  wire  uncompresser_1_0_io_decoder_ready; // @[B4Processor.scala 51:45]
  wire  uncompresser_1_0_io_decoder_valid; // @[B4Processor.scala 51:45]
  wire [31:0] uncompresser_1_0_io_decoder_bits_instruction; // @[B4Processor.scala 51:45]
  wire [63:0] uncompresser_1_0_io_decoder_bits_programCounter; // @[B4Processor.scala 51:45]
  wire  uncompresser_1_0_io_decoder_bits_wasCompressed; // @[B4Processor.scala 51:45]
  wire  decoders_0_0_io_instructionFetch_ready; // @[B4Processor.scala 54:54]
  wire  decoders_0_0_io_instructionFetch_valid; // @[B4Processor.scala 54:54]
  wire [31:0] decoders_0_0_io_instructionFetch_bits_instruction; // @[B4Processor.scala 54:54]
  wire [63:0] decoders_0_0_io_instructionFetch_bits_programCounter; // @[B4Processor.scala 54:54]
  wire  decoders_0_0_io_instructionFetch_bits_wasCompressed; // @[B4Processor.scala 54:54]
  wire [4:0] decoders_0_0_io_reorderBuffer_source1_sourceRegister; // @[B4Processor.scala 54:54]
  wire  decoders_0_0_io_reorderBuffer_source1_matchingTag_valid; // @[B4Processor.scala 54:54]
  wire [3:0] decoders_0_0_io_reorderBuffer_source1_matchingTag_bits_id; // @[B4Processor.scala 54:54]
  wire  decoders_0_0_io_reorderBuffer_source1_value_valid; // @[B4Processor.scala 54:54]
  wire [63:0] decoders_0_0_io_reorderBuffer_source1_value_bits; // @[B4Processor.scala 54:54]
  wire [4:0] decoders_0_0_io_reorderBuffer_source2_sourceRegister; // @[B4Processor.scala 54:54]
  wire  decoders_0_0_io_reorderBuffer_source2_matchingTag_valid; // @[B4Processor.scala 54:54]
  wire [3:0] decoders_0_0_io_reorderBuffer_source2_matchingTag_bits_id; // @[B4Processor.scala 54:54]
  wire  decoders_0_0_io_reorderBuffer_source2_value_valid; // @[B4Processor.scala 54:54]
  wire [63:0] decoders_0_0_io_reorderBuffer_source2_value_bits; // @[B4Processor.scala 54:54]
  wire [4:0] decoders_0_0_io_reorderBuffer_destination_destinationRegister; // @[B4Processor.scala 54:54]
  wire [3:0] decoders_0_0_io_reorderBuffer_destination_destinationTag_id; // @[B4Processor.scala 54:54]
  wire  decoders_0_0_io_reorderBuffer_destination_storeSign; // @[B4Processor.scala 54:54]
  wire  decoders_0_0_io_reorderBuffer_ready; // @[B4Processor.scala 54:54]
  wire  decoders_0_0_io_reorderBuffer_valid; // @[B4Processor.scala 54:54]
  wire  decoders_0_0_io_outputCollector_outputs_valid; // @[B4Processor.scala 54:54]
  wire  decoders_0_0_io_outputCollector_outputs_bits_resultType; // @[B4Processor.scala 54:54]
  wire [63:0] decoders_0_0_io_outputCollector_outputs_bits_value; // @[B4Processor.scala 54:54]
  wire  decoders_0_0_io_outputCollector_outputs_bits_tag_threadId; // @[B4Processor.scala 54:54]
  wire [3:0] decoders_0_0_io_outputCollector_outputs_bits_tag_id; // @[B4Processor.scala 54:54]
  wire [4:0] decoders_0_0_io_registerFile_sourceRegister1; // @[B4Processor.scala 54:54]
  wire [4:0] decoders_0_0_io_registerFile_sourceRegister2; // @[B4Processor.scala 54:54]
  wire [63:0] decoders_0_0_io_registerFile_value1; // @[B4Processor.scala 54:54]
  wire [63:0] decoders_0_0_io_registerFile_value2; // @[B4Processor.scala 54:54]
  wire  decoders_0_0_io_reservationStation_ready; // @[B4Processor.scala 54:54]
  wire [6:0] decoders_0_0_io_reservationStation_entry_opcode; // @[B4Processor.scala 54:54]
  wire [2:0] decoders_0_0_io_reservationStation_entry_function3; // @[B4Processor.scala 54:54]
  wire [11:0] decoders_0_0_io_reservationStation_entry_immediateOrFunction7; // @[B4Processor.scala 54:54]
  wire  decoders_0_0_io_reservationStation_entry_sourceTag1_threadId; // @[B4Processor.scala 54:54]
  wire [3:0] decoders_0_0_io_reservationStation_entry_sourceTag1_id; // @[B4Processor.scala 54:54]
  wire  decoders_0_0_io_reservationStation_entry_ready1; // @[B4Processor.scala 54:54]
  wire [63:0] decoders_0_0_io_reservationStation_entry_value1; // @[B4Processor.scala 54:54]
  wire  decoders_0_0_io_reservationStation_entry_sourceTag2_threadId; // @[B4Processor.scala 54:54]
  wire [3:0] decoders_0_0_io_reservationStation_entry_sourceTag2_id; // @[B4Processor.scala 54:54]
  wire  decoders_0_0_io_reservationStation_entry_ready2; // @[B4Processor.scala 54:54]
  wire [63:0] decoders_0_0_io_reservationStation_entry_value2; // @[B4Processor.scala 54:54]
  wire  decoders_0_0_io_reservationStation_entry_destinationTag_threadId; // @[B4Processor.scala 54:54]
  wire [3:0] decoders_0_0_io_reservationStation_entry_destinationTag_id; // @[B4Processor.scala 54:54]
  wire  decoders_0_0_io_reservationStation_entry_wasCompressed; // @[B4Processor.scala 54:54]
  wire  decoders_0_0_io_reservationStation_entry_valid; // @[B4Processor.scala 54:54]
  wire  decoders_0_0_io_loadStoreQueue_ready; // @[B4Processor.scala 54:54]
  wire  decoders_0_0_io_loadStoreQueue_valid; // @[B4Processor.scala 54:54]
  wire  decoders_0_0_io_loadStoreQueue_bits_accessInfo_accessType; // @[B4Processor.scala 54:54]
  wire  decoders_0_0_io_loadStoreQueue_bits_accessInfo_signed; // @[B4Processor.scala 54:54]
  wire [1:0] decoders_0_0_io_loadStoreQueue_bits_accessInfo_accessWidth; // @[B4Processor.scala 54:54]
  wire  decoders_0_0_io_loadStoreQueue_bits_addressAndLoadResultTag_threadId; // @[B4Processor.scala 54:54]
  wire [3:0] decoders_0_0_io_loadStoreQueue_bits_addressAndLoadResultTag_id; // @[B4Processor.scala 54:54]
  wire [63:0] decoders_0_0_io_loadStoreQueue_bits_address; // @[B4Processor.scala 54:54]
  wire  decoders_0_0_io_loadStoreQueue_bits_addressValid; // @[B4Processor.scala 54:54]
  wire  decoders_0_0_io_loadStoreQueue_bits_storeDataTag_threadId; // @[B4Processor.scala 54:54]
  wire [3:0] decoders_0_0_io_loadStoreQueue_bits_storeDataTag_id; // @[B4Processor.scala 54:54]
  wire [63:0] decoders_0_0_io_loadStoreQueue_bits_storeData; // @[B4Processor.scala 54:54]
  wire  decoders_0_0_io_loadStoreQueue_bits_storeDataValid; // @[B4Processor.scala 54:54]
  wire  decoders_0_0_io_csr_ready; // @[B4Processor.scala 54:54]
  wire  decoders_0_0_io_csr_valid; // @[B4Processor.scala 54:54]
  wire  decoders_0_0_io_csr_bits_sourceTag_threadId; // @[B4Processor.scala 54:54]
  wire [3:0] decoders_0_0_io_csr_bits_sourceTag_id; // @[B4Processor.scala 54:54]
  wire [3:0] decoders_0_0_io_csr_bits_destinationTag_id; // @[B4Processor.scala 54:54]
  wire [63:0] decoders_0_0_io_csr_bits_value; // @[B4Processor.scala 54:54]
  wire  decoders_0_0_io_csr_bits_ready; // @[B4Processor.scala 54:54]
  wire [11:0] decoders_0_0_io_csr_bits_address; // @[B4Processor.scala 54:54]
  wire [1:0] decoders_0_0_io_csr_bits_csrAccessType; // @[B4Processor.scala 54:54]
  wire  decoders_1_0_io_instructionFetch_ready; // @[B4Processor.scala 54:54]
  wire  decoders_1_0_io_instructionFetch_valid; // @[B4Processor.scala 54:54]
  wire [31:0] decoders_1_0_io_instructionFetch_bits_instruction; // @[B4Processor.scala 54:54]
  wire [63:0] decoders_1_0_io_instructionFetch_bits_programCounter; // @[B4Processor.scala 54:54]
  wire  decoders_1_0_io_instructionFetch_bits_wasCompressed; // @[B4Processor.scala 54:54]
  wire [4:0] decoders_1_0_io_reorderBuffer_source1_sourceRegister; // @[B4Processor.scala 54:54]
  wire  decoders_1_0_io_reorderBuffer_source1_matchingTag_valid; // @[B4Processor.scala 54:54]
  wire [3:0] decoders_1_0_io_reorderBuffer_source1_matchingTag_bits_id; // @[B4Processor.scala 54:54]
  wire  decoders_1_0_io_reorderBuffer_source1_value_valid; // @[B4Processor.scala 54:54]
  wire [63:0] decoders_1_0_io_reorderBuffer_source1_value_bits; // @[B4Processor.scala 54:54]
  wire [4:0] decoders_1_0_io_reorderBuffer_source2_sourceRegister; // @[B4Processor.scala 54:54]
  wire  decoders_1_0_io_reorderBuffer_source2_matchingTag_valid; // @[B4Processor.scala 54:54]
  wire [3:0] decoders_1_0_io_reorderBuffer_source2_matchingTag_bits_id; // @[B4Processor.scala 54:54]
  wire  decoders_1_0_io_reorderBuffer_source2_value_valid; // @[B4Processor.scala 54:54]
  wire [63:0] decoders_1_0_io_reorderBuffer_source2_value_bits; // @[B4Processor.scala 54:54]
  wire [4:0] decoders_1_0_io_reorderBuffer_destination_destinationRegister; // @[B4Processor.scala 54:54]
  wire [3:0] decoders_1_0_io_reorderBuffer_destination_destinationTag_id; // @[B4Processor.scala 54:54]
  wire  decoders_1_0_io_reorderBuffer_destination_storeSign; // @[B4Processor.scala 54:54]
  wire  decoders_1_0_io_reorderBuffer_ready; // @[B4Processor.scala 54:54]
  wire  decoders_1_0_io_reorderBuffer_valid; // @[B4Processor.scala 54:54]
  wire  decoders_1_0_io_outputCollector_outputs_valid; // @[B4Processor.scala 54:54]
  wire  decoders_1_0_io_outputCollector_outputs_bits_resultType; // @[B4Processor.scala 54:54]
  wire [63:0] decoders_1_0_io_outputCollector_outputs_bits_value; // @[B4Processor.scala 54:54]
  wire  decoders_1_0_io_outputCollector_outputs_bits_tag_threadId; // @[B4Processor.scala 54:54]
  wire [3:0] decoders_1_0_io_outputCollector_outputs_bits_tag_id; // @[B4Processor.scala 54:54]
  wire [4:0] decoders_1_0_io_registerFile_sourceRegister1; // @[B4Processor.scala 54:54]
  wire [4:0] decoders_1_0_io_registerFile_sourceRegister2; // @[B4Processor.scala 54:54]
  wire [63:0] decoders_1_0_io_registerFile_value1; // @[B4Processor.scala 54:54]
  wire [63:0] decoders_1_0_io_registerFile_value2; // @[B4Processor.scala 54:54]
  wire  decoders_1_0_io_reservationStation_ready; // @[B4Processor.scala 54:54]
  wire [6:0] decoders_1_0_io_reservationStation_entry_opcode; // @[B4Processor.scala 54:54]
  wire [2:0] decoders_1_0_io_reservationStation_entry_function3; // @[B4Processor.scala 54:54]
  wire [11:0] decoders_1_0_io_reservationStation_entry_immediateOrFunction7; // @[B4Processor.scala 54:54]
  wire  decoders_1_0_io_reservationStation_entry_sourceTag1_threadId; // @[B4Processor.scala 54:54]
  wire [3:0] decoders_1_0_io_reservationStation_entry_sourceTag1_id; // @[B4Processor.scala 54:54]
  wire  decoders_1_0_io_reservationStation_entry_ready1; // @[B4Processor.scala 54:54]
  wire [63:0] decoders_1_0_io_reservationStation_entry_value1; // @[B4Processor.scala 54:54]
  wire  decoders_1_0_io_reservationStation_entry_sourceTag2_threadId; // @[B4Processor.scala 54:54]
  wire [3:0] decoders_1_0_io_reservationStation_entry_sourceTag2_id; // @[B4Processor.scala 54:54]
  wire  decoders_1_0_io_reservationStation_entry_ready2; // @[B4Processor.scala 54:54]
  wire [63:0] decoders_1_0_io_reservationStation_entry_value2; // @[B4Processor.scala 54:54]
  wire  decoders_1_0_io_reservationStation_entry_destinationTag_threadId; // @[B4Processor.scala 54:54]
  wire [3:0] decoders_1_0_io_reservationStation_entry_destinationTag_id; // @[B4Processor.scala 54:54]
  wire  decoders_1_0_io_reservationStation_entry_wasCompressed; // @[B4Processor.scala 54:54]
  wire  decoders_1_0_io_reservationStation_entry_valid; // @[B4Processor.scala 54:54]
  wire  decoders_1_0_io_loadStoreQueue_ready; // @[B4Processor.scala 54:54]
  wire  decoders_1_0_io_loadStoreQueue_valid; // @[B4Processor.scala 54:54]
  wire  decoders_1_0_io_loadStoreQueue_bits_accessInfo_accessType; // @[B4Processor.scala 54:54]
  wire  decoders_1_0_io_loadStoreQueue_bits_accessInfo_signed; // @[B4Processor.scala 54:54]
  wire [1:0] decoders_1_0_io_loadStoreQueue_bits_accessInfo_accessWidth; // @[B4Processor.scala 54:54]
  wire  decoders_1_0_io_loadStoreQueue_bits_addressAndLoadResultTag_threadId; // @[B4Processor.scala 54:54]
  wire [3:0] decoders_1_0_io_loadStoreQueue_bits_addressAndLoadResultTag_id; // @[B4Processor.scala 54:54]
  wire [63:0] decoders_1_0_io_loadStoreQueue_bits_address; // @[B4Processor.scala 54:54]
  wire  decoders_1_0_io_loadStoreQueue_bits_addressValid; // @[B4Processor.scala 54:54]
  wire  decoders_1_0_io_loadStoreQueue_bits_storeDataTag_threadId; // @[B4Processor.scala 54:54]
  wire [3:0] decoders_1_0_io_loadStoreQueue_bits_storeDataTag_id; // @[B4Processor.scala 54:54]
  wire [63:0] decoders_1_0_io_loadStoreQueue_bits_storeData; // @[B4Processor.scala 54:54]
  wire  decoders_1_0_io_loadStoreQueue_bits_storeDataValid; // @[B4Processor.scala 54:54]
  wire  decoders_1_0_io_csr_ready; // @[B4Processor.scala 54:54]
  wire  decoders_1_0_io_csr_valid; // @[B4Processor.scala 54:54]
  wire  decoders_1_0_io_csr_bits_sourceTag_threadId; // @[B4Processor.scala 54:54]
  wire [3:0] decoders_1_0_io_csr_bits_sourceTag_id; // @[B4Processor.scala 54:54]
  wire [3:0] decoders_1_0_io_csr_bits_destinationTag_id; // @[B4Processor.scala 54:54]
  wire [63:0] decoders_1_0_io_csr_bits_value; // @[B4Processor.scala 54:54]
  wire  decoders_1_0_io_csr_bits_ready; // @[B4Processor.scala 54:54]
  wire [11:0] decoders_1_0_io_csr_bits_address; // @[B4Processor.scala 54:54]
  wire [1:0] decoders_1_0_io_csr_bits_csrAccessType; // @[B4Processor.scala 54:54]
  wire  reservationStation_clock; // @[B4Processor.scala 56:42]
  wire  reservationStation_reset; // @[B4Processor.scala 56:42]
  wire  reservationStation_io_collectedOutput_0_outputs_valid; // @[B4Processor.scala 56:42]
  wire  reservationStation_io_collectedOutput_0_outputs_bits_resultType; // @[B4Processor.scala 56:42]
  wire [63:0] reservationStation_io_collectedOutput_0_outputs_bits_value; // @[B4Processor.scala 56:42]
  wire  reservationStation_io_collectedOutput_0_outputs_bits_tag_threadId; // @[B4Processor.scala 56:42]
  wire [3:0] reservationStation_io_collectedOutput_0_outputs_bits_tag_id; // @[B4Processor.scala 56:42]
  wire  reservationStation_io_collectedOutput_1_outputs_valid; // @[B4Processor.scala 56:42]
  wire  reservationStation_io_collectedOutput_1_outputs_bits_resultType; // @[B4Processor.scala 56:42]
  wire [63:0] reservationStation_io_collectedOutput_1_outputs_bits_value; // @[B4Processor.scala 56:42]
  wire  reservationStation_io_collectedOutput_1_outputs_bits_tag_threadId; // @[B4Processor.scala 56:42]
  wire [3:0] reservationStation_io_collectedOutput_1_outputs_bits_tag_id; // @[B4Processor.scala 56:42]
  wire  reservationStation_io_executor_0_ready; // @[B4Processor.scala 56:42]
  wire  reservationStation_io_executor_0_valid; // @[B4Processor.scala 56:42]
  wire  reservationStation_io_executor_0_bits_destinationTag_threadId; // @[B4Processor.scala 56:42]
  wire [3:0] reservationStation_io_executor_0_bits_destinationTag_id; // @[B4Processor.scala 56:42]
  wire [63:0] reservationStation_io_executor_0_bits_value1; // @[B4Processor.scala 56:42]
  wire [63:0] reservationStation_io_executor_0_bits_value2; // @[B4Processor.scala 56:42]
  wire [2:0] reservationStation_io_executor_0_bits_function3; // @[B4Processor.scala 56:42]
  wire [11:0] reservationStation_io_executor_0_bits_immediateOrFunction7; // @[B4Processor.scala 56:42]
  wire [6:0] reservationStation_io_executor_0_bits_opcode; // @[B4Processor.scala 56:42]
  wire  reservationStation_io_executor_0_bits_wasCompressed; // @[B4Processor.scala 56:42]
  wire  reservationStation_io_executor_1_ready; // @[B4Processor.scala 56:42]
  wire  reservationStation_io_executor_1_valid; // @[B4Processor.scala 56:42]
  wire  reservationStation_io_executor_1_bits_destinationTag_threadId; // @[B4Processor.scala 56:42]
  wire [3:0] reservationStation_io_executor_1_bits_destinationTag_id; // @[B4Processor.scala 56:42]
  wire [63:0] reservationStation_io_executor_1_bits_value1; // @[B4Processor.scala 56:42]
  wire [63:0] reservationStation_io_executor_1_bits_value2; // @[B4Processor.scala 56:42]
  wire [2:0] reservationStation_io_executor_1_bits_function3; // @[B4Processor.scala 56:42]
  wire [11:0] reservationStation_io_executor_1_bits_immediateOrFunction7; // @[B4Processor.scala 56:42]
  wire [6:0] reservationStation_io_executor_1_bits_opcode; // @[B4Processor.scala 56:42]
  wire  reservationStation_io_executor_1_bits_wasCompressed; // @[B4Processor.scala 56:42]
  wire  reservationStation_io_decoder_0_ready; // @[B4Processor.scala 56:42]
  wire [6:0] reservationStation_io_decoder_0_entry_opcode; // @[B4Processor.scala 56:42]
  wire [2:0] reservationStation_io_decoder_0_entry_function3; // @[B4Processor.scala 56:42]
  wire [11:0] reservationStation_io_decoder_0_entry_immediateOrFunction7; // @[B4Processor.scala 56:42]
  wire  reservationStation_io_decoder_0_entry_sourceTag1_threadId; // @[B4Processor.scala 56:42]
  wire [3:0] reservationStation_io_decoder_0_entry_sourceTag1_id; // @[B4Processor.scala 56:42]
  wire  reservationStation_io_decoder_0_entry_ready1; // @[B4Processor.scala 56:42]
  wire [63:0] reservationStation_io_decoder_0_entry_value1; // @[B4Processor.scala 56:42]
  wire  reservationStation_io_decoder_0_entry_sourceTag2_threadId; // @[B4Processor.scala 56:42]
  wire [3:0] reservationStation_io_decoder_0_entry_sourceTag2_id; // @[B4Processor.scala 56:42]
  wire  reservationStation_io_decoder_0_entry_ready2; // @[B4Processor.scala 56:42]
  wire [63:0] reservationStation_io_decoder_0_entry_value2; // @[B4Processor.scala 56:42]
  wire [3:0] reservationStation_io_decoder_0_entry_destinationTag_id; // @[B4Processor.scala 56:42]
  wire  reservationStation_io_decoder_0_entry_wasCompressed; // @[B4Processor.scala 56:42]
  wire  reservationStation_io_decoder_0_entry_valid; // @[B4Processor.scala 56:42]
  wire  reservationStation_io_decoder_1_ready; // @[B4Processor.scala 56:42]
  wire [6:0] reservationStation_io_decoder_1_entry_opcode; // @[B4Processor.scala 56:42]
  wire [2:0] reservationStation_io_decoder_1_entry_function3; // @[B4Processor.scala 56:42]
  wire [11:0] reservationStation_io_decoder_1_entry_immediateOrFunction7; // @[B4Processor.scala 56:42]
  wire  reservationStation_io_decoder_1_entry_sourceTag1_threadId; // @[B4Processor.scala 56:42]
  wire [3:0] reservationStation_io_decoder_1_entry_sourceTag1_id; // @[B4Processor.scala 56:42]
  wire  reservationStation_io_decoder_1_entry_ready1; // @[B4Processor.scala 56:42]
  wire [63:0] reservationStation_io_decoder_1_entry_value1; // @[B4Processor.scala 56:42]
  wire  reservationStation_io_decoder_1_entry_sourceTag2_threadId; // @[B4Processor.scala 56:42]
  wire [3:0] reservationStation_io_decoder_1_entry_sourceTag2_id; // @[B4Processor.scala 56:42]
  wire  reservationStation_io_decoder_1_entry_ready2; // @[B4Processor.scala 56:42]
  wire [63:0] reservationStation_io_decoder_1_entry_value2; // @[B4Processor.scala 56:42]
  wire [3:0] reservationStation_io_decoder_1_entry_destinationTag_id; // @[B4Processor.scala 56:42]
  wire  reservationStation_io_decoder_1_entry_wasCompressed; // @[B4Processor.scala 56:42]
  wire  reservationStation_io_decoder_1_entry_valid; // @[B4Processor.scala 56:42]
  wire  executors_0_io_reservationStation_ready; // @[B4Processor.scala 57:60]
  wire  executors_0_io_reservationStation_valid; // @[B4Processor.scala 57:60]
  wire  executors_0_io_reservationStation_bits_destinationTag_threadId; // @[B4Processor.scala 57:60]
  wire [3:0] executors_0_io_reservationStation_bits_destinationTag_id; // @[B4Processor.scala 57:60]
  wire [63:0] executors_0_io_reservationStation_bits_value1; // @[B4Processor.scala 57:60]
  wire [63:0] executors_0_io_reservationStation_bits_value2; // @[B4Processor.scala 57:60]
  wire [2:0] executors_0_io_reservationStation_bits_function3; // @[B4Processor.scala 57:60]
  wire [11:0] executors_0_io_reservationStation_bits_immediateOrFunction7; // @[B4Processor.scala 57:60]
  wire [6:0] executors_0_io_reservationStation_bits_opcode; // @[B4Processor.scala 57:60]
  wire  executors_0_io_reservationStation_bits_wasCompressed; // @[B4Processor.scala 57:60]
  wire  executors_0_io_out_ready; // @[B4Processor.scala 57:60]
  wire  executors_0_io_out_valid; // @[B4Processor.scala 57:60]
  wire  executors_0_io_out_bits_resultType; // @[B4Processor.scala 57:60]
  wire [63:0] executors_0_io_out_bits_value; // @[B4Processor.scala 57:60]
  wire  executors_0_io_out_bits_tag_threadId; // @[B4Processor.scala 57:60]
  wire [3:0] executors_0_io_out_bits_tag_id; // @[B4Processor.scala 57:60]
  wire  executors_0_io_fetch_ready; // @[B4Processor.scala 57:60]
  wire  executors_0_io_fetch_valid; // @[B4Processor.scala 57:60]
  wire  executors_0_io_fetch_bits_threadId; // @[B4Processor.scala 57:60]
  wire [63:0] executors_0_io_fetch_bits_programCounterOffset; // @[B4Processor.scala 57:60]
  wire  executors_1_io_reservationStation_ready; // @[B4Processor.scala 57:60]
  wire  executors_1_io_reservationStation_valid; // @[B4Processor.scala 57:60]
  wire  executors_1_io_reservationStation_bits_destinationTag_threadId; // @[B4Processor.scala 57:60]
  wire [3:0] executors_1_io_reservationStation_bits_destinationTag_id; // @[B4Processor.scala 57:60]
  wire [63:0] executors_1_io_reservationStation_bits_value1; // @[B4Processor.scala 57:60]
  wire [63:0] executors_1_io_reservationStation_bits_value2; // @[B4Processor.scala 57:60]
  wire [2:0] executors_1_io_reservationStation_bits_function3; // @[B4Processor.scala 57:60]
  wire [11:0] executors_1_io_reservationStation_bits_immediateOrFunction7; // @[B4Processor.scala 57:60]
  wire [6:0] executors_1_io_reservationStation_bits_opcode; // @[B4Processor.scala 57:60]
  wire  executors_1_io_reservationStation_bits_wasCompressed; // @[B4Processor.scala 57:60]
  wire  executors_1_io_out_ready; // @[B4Processor.scala 57:60]
  wire  executors_1_io_out_valid; // @[B4Processor.scala 57:60]
  wire  executors_1_io_out_bits_resultType; // @[B4Processor.scala 57:60]
  wire [63:0] executors_1_io_out_bits_value; // @[B4Processor.scala 57:60]
  wire  executors_1_io_out_bits_tag_threadId; // @[B4Processor.scala 57:60]
  wire [3:0] executors_1_io_out_bits_tag_id; // @[B4Processor.scala 57:60]
  wire  executors_1_io_fetch_ready; // @[B4Processor.scala 57:60]
  wire  executors_1_io_fetch_valid; // @[B4Processor.scala 57:60]
  wire  executors_1_io_fetch_bits_threadId; // @[B4Processor.scala 57:60]
  wire [63:0] executors_1_io_fetch_bits_programCounterOffset; // @[B4Processor.scala 57:60]
  wire  externalMemoryInterface_clock; // @[B4Processor.scala 59:47]
  wire  externalMemoryInterface_reset; // @[B4Processor.scala 59:47]
  wire  externalMemoryInterface_io_dataWriteRequests_ready; // @[B4Processor.scala 59:47]
  wire  externalMemoryInterface_io_dataWriteRequests_valid; // @[B4Processor.scala 59:47]
  wire [63:0] externalMemoryInterface_io_dataWriteRequests_bits_address; // @[B4Processor.scala 59:47]
  wire [63:0] externalMemoryInterface_io_dataWriteRequests_bits_data; // @[B4Processor.scala 59:47]
  wire [7:0] externalMemoryInterface_io_dataWriteRequests_bits_mask; // @[B4Processor.scala 59:47]
  wire  externalMemoryInterface_io_dataReadRequests_ready; // @[B4Processor.scala 59:47]
  wire  externalMemoryInterface_io_dataReadRequests_valid; // @[B4Processor.scala 59:47]
  wire [63:0] externalMemoryInterface_io_dataReadRequests_bits_address; // @[B4Processor.scala 59:47]
  wire [1:0] externalMemoryInterface_io_dataReadRequests_bits_size; // @[B4Processor.scala 59:47]
  wire  externalMemoryInterface_io_dataReadRequests_bits_signed; // @[B4Processor.scala 59:47]
  wire  externalMemoryInterface_io_dataReadRequests_bits_outputTag_threadId; // @[B4Processor.scala 59:47]
  wire [3:0] externalMemoryInterface_io_dataReadRequests_bits_outputTag_id; // @[B4Processor.scala 59:47]
  wire  externalMemoryInterface_io_instructionFetchRequest_0_ready; // @[B4Processor.scala 59:47]
  wire  externalMemoryInterface_io_instructionFetchRequest_0_valid; // @[B4Processor.scala 59:47]
  wire [63:0] externalMemoryInterface_io_instructionFetchRequest_0_bits_address; // @[B4Processor.scala 59:47]
  wire  externalMemoryInterface_io_instructionFetchRequest_1_ready; // @[B4Processor.scala 59:47]
  wire  externalMemoryInterface_io_instructionFetchRequest_1_valid; // @[B4Processor.scala 59:47]
  wire [63:0] externalMemoryInterface_io_instructionFetchRequest_1_bits_address; // @[B4Processor.scala 59:47]
  wire  externalMemoryInterface_io_dataReadOut_ready; // @[B4Processor.scala 59:47]
  wire  externalMemoryInterface_io_dataReadOut_valid; // @[B4Processor.scala 59:47]
  wire [63:0] externalMemoryInterface_io_dataReadOut_bits_value; // @[B4Processor.scala 59:47]
  wire  externalMemoryInterface_io_dataReadOut_bits_isError; // @[B4Processor.scala 59:47]
  wire  externalMemoryInterface_io_dataReadOut_bits_tag_threadId; // @[B4Processor.scala 59:47]
  wire [3:0] externalMemoryInterface_io_dataReadOut_bits_tag_id; // @[B4Processor.scala 59:47]
  wire  externalMemoryInterface_io_instructionOut_0_valid; // @[B4Processor.scala 59:47]
  wire [63:0] externalMemoryInterface_io_instructionOut_0_bits_inner; // @[B4Processor.scala 59:47]
  wire  externalMemoryInterface_io_instructionOut_1_valid; // @[B4Processor.scala 59:47]
  wire [63:0] externalMemoryInterface_io_instructionOut_1_bits_inner; // @[B4Processor.scala 59:47]
  wire  externalMemoryInterface_io_coordinator_writeAddress_ready; // @[B4Processor.scala 59:47]
  wire  externalMemoryInterface_io_coordinator_writeAddress_valid; // @[B4Processor.scala 59:47]
  wire [63:0] externalMemoryInterface_io_coordinator_writeAddress_bits_ADDR; // @[B4Processor.scala 59:47]
  wire [3:0] externalMemoryInterface_io_coordinator_writeAddress_bits_CACHE; // @[B4Processor.scala 59:47]
  wire  externalMemoryInterface_io_coordinator_write_ready; // @[B4Processor.scala 59:47]
  wire  externalMemoryInterface_io_coordinator_write_valid; // @[B4Processor.scala 59:47]
  wire [63:0] externalMemoryInterface_io_coordinator_write_bits_DATA; // @[B4Processor.scala 59:47]
  wire [7:0] externalMemoryInterface_io_coordinator_write_bits_STRB; // @[B4Processor.scala 59:47]
  wire  externalMemoryInterface_io_coordinator_write_bits_LAST; // @[B4Processor.scala 59:47]
  wire  externalMemoryInterface_io_coordinator_writeResponse_ready; // @[B4Processor.scala 59:47]
  wire  externalMemoryInterface_io_coordinator_writeResponse_valid; // @[B4Processor.scala 59:47]
  wire  externalMemoryInterface_io_coordinator_readAddress_ready; // @[B4Processor.scala 59:47]
  wire  externalMemoryInterface_io_coordinator_readAddress_valid; // @[B4Processor.scala 59:47]
  wire [63:0] externalMemoryInterface_io_coordinator_readAddress_bits_ADDR; // @[B4Processor.scala 59:47]
  wire [7:0] externalMemoryInterface_io_coordinator_readAddress_bits_LEN; // @[B4Processor.scala 59:47]
  wire [3:0] externalMemoryInterface_io_coordinator_readAddress_bits_CACHE; // @[B4Processor.scala 59:47]
  wire  externalMemoryInterface_io_coordinator_read_ready; // @[B4Processor.scala 59:47]
  wire  externalMemoryInterface_io_coordinator_read_valid; // @[B4Processor.scala 59:47]
  wire [63:0] externalMemoryInterface_io_coordinator_read_bits_DATA; // @[B4Processor.scala 59:47]
  wire [1:0] externalMemoryInterface_io_coordinator_read_bits_RESP; // @[B4Processor.scala 59:47]
  wire  csrReservationStation_0_clock; // @[B4Processor.scala 62:36]
  wire  csrReservationStation_0_reset; // @[B4Processor.scala 62:36]
  wire  csrReservationStation_0_io_decoderInput_0_ready; // @[B4Processor.scala 62:36]
  wire  csrReservationStation_0_io_decoderInput_0_valid; // @[B4Processor.scala 62:36]
  wire  csrReservationStation_0_io_decoderInput_0_bits_sourceTag_threadId; // @[B4Processor.scala 62:36]
  wire [3:0] csrReservationStation_0_io_decoderInput_0_bits_sourceTag_id; // @[B4Processor.scala 62:36]
  wire  csrReservationStation_0_io_decoderInput_0_bits_destinationTag_threadId; // @[B4Processor.scala 62:36]
  wire [3:0] csrReservationStation_0_io_decoderInput_0_bits_destinationTag_id; // @[B4Processor.scala 62:36]
  wire [63:0] csrReservationStation_0_io_decoderInput_0_bits_value; // @[B4Processor.scala 62:36]
  wire  csrReservationStation_0_io_decoderInput_0_bits_ready; // @[B4Processor.scala 62:36]
  wire [11:0] csrReservationStation_0_io_decoderInput_0_bits_address; // @[B4Processor.scala 62:36]
  wire [1:0] csrReservationStation_0_io_decoderInput_0_bits_csrAccessType; // @[B4Processor.scala 62:36]
  wire  csrReservationStation_0_io_toCSR_ready; // @[B4Processor.scala 62:36]
  wire  csrReservationStation_0_io_toCSR_valid; // @[B4Processor.scala 62:36]
  wire [11:0] csrReservationStation_0_io_toCSR_bits_address; // @[B4Processor.scala 62:36]
  wire [63:0] csrReservationStation_0_io_toCSR_bits_value; // @[B4Processor.scala 62:36]
  wire  csrReservationStation_0_io_toCSR_bits_destinationTag_threadId; // @[B4Processor.scala 62:36]
  wire [3:0] csrReservationStation_0_io_toCSR_bits_destinationTag_id; // @[B4Processor.scala 62:36]
  wire [1:0] csrReservationStation_0_io_toCSR_bits_csrAccessType; // @[B4Processor.scala 62:36]
  wire  csrReservationStation_0_io_output_outputs_valid; // @[B4Processor.scala 62:36]
  wire [63:0] csrReservationStation_0_io_output_outputs_bits_value; // @[B4Processor.scala 62:36]
  wire  csrReservationStation_0_io_output_outputs_bits_tag_threadId; // @[B4Processor.scala 62:36]
  wire [3:0] csrReservationStation_0_io_output_outputs_bits_tag_id; // @[B4Processor.scala 62:36]
  wire  csrReservationStation_0_io_empty; // @[B4Processor.scala 62:36]
  wire  csrReservationStation_1_clock; // @[B4Processor.scala 62:36]
  wire  csrReservationStation_1_reset; // @[B4Processor.scala 62:36]
  wire  csrReservationStation_1_io_decoderInput_0_ready; // @[B4Processor.scala 62:36]
  wire  csrReservationStation_1_io_decoderInput_0_valid; // @[B4Processor.scala 62:36]
  wire  csrReservationStation_1_io_decoderInput_0_bits_sourceTag_threadId; // @[B4Processor.scala 62:36]
  wire [3:0] csrReservationStation_1_io_decoderInput_0_bits_sourceTag_id; // @[B4Processor.scala 62:36]
  wire  csrReservationStation_1_io_decoderInput_0_bits_destinationTag_threadId; // @[B4Processor.scala 62:36]
  wire [3:0] csrReservationStation_1_io_decoderInput_0_bits_destinationTag_id; // @[B4Processor.scala 62:36]
  wire [63:0] csrReservationStation_1_io_decoderInput_0_bits_value; // @[B4Processor.scala 62:36]
  wire  csrReservationStation_1_io_decoderInput_0_bits_ready; // @[B4Processor.scala 62:36]
  wire [11:0] csrReservationStation_1_io_decoderInput_0_bits_address; // @[B4Processor.scala 62:36]
  wire [1:0] csrReservationStation_1_io_decoderInput_0_bits_csrAccessType; // @[B4Processor.scala 62:36]
  wire  csrReservationStation_1_io_toCSR_ready; // @[B4Processor.scala 62:36]
  wire  csrReservationStation_1_io_toCSR_valid; // @[B4Processor.scala 62:36]
  wire [11:0] csrReservationStation_1_io_toCSR_bits_address; // @[B4Processor.scala 62:36]
  wire [63:0] csrReservationStation_1_io_toCSR_bits_value; // @[B4Processor.scala 62:36]
  wire  csrReservationStation_1_io_toCSR_bits_destinationTag_threadId; // @[B4Processor.scala 62:36]
  wire [3:0] csrReservationStation_1_io_toCSR_bits_destinationTag_id; // @[B4Processor.scala 62:36]
  wire [1:0] csrReservationStation_1_io_toCSR_bits_csrAccessType; // @[B4Processor.scala 62:36]
  wire  csrReservationStation_1_io_output_outputs_valid; // @[B4Processor.scala 62:36]
  wire [63:0] csrReservationStation_1_io_output_outputs_bits_value; // @[B4Processor.scala 62:36]
  wire  csrReservationStation_1_io_output_outputs_bits_tag_threadId; // @[B4Processor.scala 62:36]
  wire [3:0] csrReservationStation_1_io_output_outputs_bits_tag_id; // @[B4Processor.scala 62:36]
  wire  csrReservationStation_1_io_empty; // @[B4Processor.scala 62:36]
  wire  csr_0_clock; // @[B4Processor.scala 63:61]
  wire  csr_0_reset; // @[B4Processor.scala 63:61]
  wire  csr_0_io_decoderInput_ready; // @[B4Processor.scala 63:61]
  wire  csr_0_io_decoderInput_valid; // @[B4Processor.scala 63:61]
  wire [11:0] csr_0_io_decoderInput_bits_address; // @[B4Processor.scala 63:61]
  wire [63:0] csr_0_io_decoderInput_bits_value; // @[B4Processor.scala 63:61]
  wire  csr_0_io_decoderInput_bits_destinationTag_threadId; // @[B4Processor.scala 63:61]
  wire [3:0] csr_0_io_decoderInput_bits_destinationTag_id; // @[B4Processor.scala 63:61]
  wire [1:0] csr_0_io_decoderInput_bits_csrAccessType; // @[B4Processor.scala 63:61]
  wire  csr_0_io_CSROutput_ready; // @[B4Processor.scala 63:61]
  wire  csr_0_io_CSROutput_valid; // @[B4Processor.scala 63:61]
  wire [63:0] csr_0_io_CSROutput_bits_value; // @[B4Processor.scala 63:61]
  wire  csr_0_io_CSROutput_bits_isError; // @[B4Processor.scala 63:61]
  wire  csr_0_io_CSROutput_bits_tag_threadId; // @[B4Processor.scala 63:61]
  wire [3:0] csr_0_io_CSROutput_bits_tag_id; // @[B4Processor.scala 63:61]
  wire [63:0] csr_0_io_fetch_mtvec; // @[B4Processor.scala 63:61]
  wire [63:0] csr_0_io_fetch_mepc; // @[B4Processor.scala 63:61]
  wire [63:0] csr_0_io_fetch_mcause; // @[B4Processor.scala 63:61]
  wire [1:0] csr_0_io_reorderBuffer_retireCount; // @[B4Processor.scala 63:61]
  wire  csr_1_clock; // @[B4Processor.scala 63:61]
  wire  csr_1_reset; // @[B4Processor.scala 63:61]
  wire  csr_1_io_decoderInput_ready; // @[B4Processor.scala 63:61]
  wire  csr_1_io_decoderInput_valid; // @[B4Processor.scala 63:61]
  wire [11:0] csr_1_io_decoderInput_bits_address; // @[B4Processor.scala 63:61]
  wire [63:0] csr_1_io_decoderInput_bits_value; // @[B4Processor.scala 63:61]
  wire  csr_1_io_decoderInput_bits_destinationTag_threadId; // @[B4Processor.scala 63:61]
  wire [3:0] csr_1_io_decoderInput_bits_destinationTag_id; // @[B4Processor.scala 63:61]
  wire [1:0] csr_1_io_decoderInput_bits_csrAccessType; // @[B4Processor.scala 63:61]
  wire  csr_1_io_CSROutput_ready; // @[B4Processor.scala 63:61]
  wire  csr_1_io_CSROutput_valid; // @[B4Processor.scala 63:61]
  wire [63:0] csr_1_io_CSROutput_bits_value; // @[B4Processor.scala 63:61]
  wire  csr_1_io_CSROutput_bits_isError; // @[B4Processor.scala 63:61]
  wire  csr_1_io_CSROutput_bits_tag_threadId; // @[B4Processor.scala 63:61]
  wire [3:0] csr_1_io_CSROutput_bits_tag_id; // @[B4Processor.scala 63:61]
  wire [63:0] csr_1_io_fetch_mtvec; // @[B4Processor.scala 63:61]
  wire [63:0] csr_1_io_fetch_mepc; // @[B4Processor.scala 63:61]
  wire [63:0] csr_1_io_fetch_mcause; // @[B4Processor.scala 63:61]
  wire [1:0] csr_1_io_reorderBuffer_retireCount; // @[B4Processor.scala 63:61]
  InstructionMemoryCache instructionCache_0 ( // @[B4Processor.scala 35:45]
    .clock(instructionCache_0_clock),
    .reset(instructionCache_0_reset),
    .io_fetch_0_address_valid(instructionCache_0_io_fetch_0_address_valid),
    .io_fetch_0_address_bits(instructionCache_0_io_fetch_0_address_bits),
    .io_fetch_0_output_valid(instructionCache_0_io_fetch_0_output_valid),
    .io_fetch_0_output_bits(instructionCache_0_io_fetch_0_output_bits),
    .io_memory_request_ready(instructionCache_0_io_memory_request_ready),
    .io_memory_request_valid(instructionCache_0_io_memory_request_valid),
    .io_memory_request_bits_address(instructionCache_0_io_memory_request_bits_address),
    .io_memory_response_valid(instructionCache_0_io_memory_response_valid),
    .io_memory_response_bits_inner(instructionCache_0_io_memory_response_bits_inner)
  );
  InstructionMemoryCache_1 instructionCache_1 ( // @[B4Processor.scala 35:45]
    .clock(instructionCache_1_clock),
    .reset(instructionCache_1_reset),
    .io_fetch_0_address_valid(instructionCache_1_io_fetch_0_address_valid),
    .io_fetch_0_address_bits(instructionCache_1_io_fetch_0_address_bits),
    .io_fetch_0_output_valid(instructionCache_1_io_fetch_0_output_valid),
    .io_fetch_0_output_bits(instructionCache_1_io_fetch_0_output_bits),
    .io_memory_request_ready(instructionCache_1_io_memory_request_ready),
    .io_memory_request_valid(instructionCache_1_io_memory_request_valid),
    .io_memory_request_bits_address(instructionCache_1_io_memory_request_bits_address),
    .io_memory_response_valid(instructionCache_1_io_memory_response_valid),
    .io_memory_response_bits_inner(instructionCache_1_io_memory_response_bits_inner)
  );
  Fetch fetch_0 ( // @[B4Processor.scala 36:63]
    .clock(fetch_0_clock),
    .reset(fetch_0_reset),
    .io_cache_0_address_valid(fetch_0_io_cache_0_address_valid),
    .io_cache_0_address_bits(fetch_0_io_cache_0_address_bits),
    .io_cache_0_output_valid(fetch_0_io_cache_0_output_valid),
    .io_cache_0_output_bits(fetch_0_io_cache_0_output_bits),
    .io_reorderBufferEmpty(fetch_0_io_reorderBufferEmpty),
    .io_loadStoreQueueEmpty(fetch_0_io_loadStoreQueueEmpty),
    .io_collectedBranchAddresses_addresses_valid(fetch_0_io_collectedBranchAddresses_addresses_valid),
    .io_collectedBranchAddresses_addresses_bits_threadId(fetch_0_io_collectedBranchAddresses_addresses_bits_threadId),
    .io_collectedBranchAddresses_addresses_bits_programCounterOffset(
      fetch_0_io_collectedBranchAddresses_addresses_bits_programCounterOffset),
    .io_fetchBuffer_toBuffer_0_ready(fetch_0_io_fetchBuffer_toBuffer_0_ready),
    .io_fetchBuffer_toBuffer_0_valid(fetch_0_io_fetchBuffer_toBuffer_0_valid),
    .io_fetchBuffer_toBuffer_0_bits_instruction(fetch_0_io_fetchBuffer_toBuffer_0_bits_instruction),
    .io_fetchBuffer_toBuffer_0_bits_programCounter(fetch_0_io_fetchBuffer_toBuffer_0_bits_programCounter),
    .io_fetchBuffer_empty(fetch_0_io_fetchBuffer_empty),
    .io_csr_mtvec(fetch_0_io_csr_mtvec),
    .io_csr_mepc(fetch_0_io_csr_mepc),
    .io_csr_mcause(fetch_0_io_csr_mcause),
    .io_csrReservationStationEmpty(fetch_0_io_csrReservationStationEmpty),
    .io_isError(fetch_0_io_isError)
  );
  Fetch_1 fetch_1 ( // @[B4Processor.scala 36:63]
    .clock(fetch_1_clock),
    .reset(fetch_1_reset),
    .io_cache_0_address_valid(fetch_1_io_cache_0_address_valid),
    .io_cache_0_address_bits(fetch_1_io_cache_0_address_bits),
    .io_cache_0_output_valid(fetch_1_io_cache_0_output_valid),
    .io_cache_0_output_bits(fetch_1_io_cache_0_output_bits),
    .io_reorderBufferEmpty(fetch_1_io_reorderBufferEmpty),
    .io_loadStoreQueueEmpty(fetch_1_io_loadStoreQueueEmpty),
    .io_collectedBranchAddresses_addresses_valid(fetch_1_io_collectedBranchAddresses_addresses_valid),
    .io_collectedBranchAddresses_addresses_bits_threadId(fetch_1_io_collectedBranchAddresses_addresses_bits_threadId),
    .io_collectedBranchAddresses_addresses_bits_programCounterOffset(
      fetch_1_io_collectedBranchAddresses_addresses_bits_programCounterOffset),
    .io_fetchBuffer_toBuffer_0_ready(fetch_1_io_fetchBuffer_toBuffer_0_ready),
    .io_fetchBuffer_toBuffer_0_valid(fetch_1_io_fetchBuffer_toBuffer_0_valid),
    .io_fetchBuffer_toBuffer_0_bits_instruction(fetch_1_io_fetchBuffer_toBuffer_0_bits_instruction),
    .io_fetchBuffer_toBuffer_0_bits_programCounter(fetch_1_io_fetchBuffer_toBuffer_0_bits_programCounter),
    .io_fetchBuffer_empty(fetch_1_io_fetchBuffer_empty),
    .io_csr_mtvec(fetch_1_io_csr_mtvec),
    .io_csr_mepc(fetch_1_io_csr_mepc),
    .io_csr_mcause(fetch_1_io_csr_mcause),
    .io_csrReservationStationEmpty(fetch_1_io_csrReservationStationEmpty),
    .io_isError(fetch_1_io_isError)
  );
  FetchBuffer fetchBuffer_0 ( // @[B4Processor.scala 38:45]
    .clock(fetchBuffer_0_clock),
    .reset(fetchBuffer_0_reset),
    .io_output_0_ready(fetchBuffer_0_io_output_0_ready),
    .io_output_0_valid(fetchBuffer_0_io_output_0_valid),
    .io_output_0_bits_instruction(fetchBuffer_0_io_output_0_bits_instruction),
    .io_output_0_bits_programCounter(fetchBuffer_0_io_output_0_bits_programCounter),
    .io_input_toBuffer_0_ready(fetchBuffer_0_io_input_toBuffer_0_ready),
    .io_input_toBuffer_0_valid(fetchBuffer_0_io_input_toBuffer_0_valid),
    .io_input_toBuffer_0_bits_instruction(fetchBuffer_0_io_input_toBuffer_0_bits_instruction),
    .io_input_toBuffer_0_bits_programCounter(fetchBuffer_0_io_input_toBuffer_0_bits_programCounter),
    .io_input_empty(fetchBuffer_0_io_input_empty)
  );
  FetchBuffer fetchBuffer_1 ( // @[B4Processor.scala 38:45]
    .clock(fetchBuffer_1_clock),
    .reset(fetchBuffer_1_reset),
    .io_output_0_ready(fetchBuffer_1_io_output_0_ready),
    .io_output_0_valid(fetchBuffer_1_io_output_0_valid),
    .io_output_0_bits_instruction(fetchBuffer_1_io_output_0_bits_instruction),
    .io_output_0_bits_programCounter(fetchBuffer_1_io_output_0_bits_programCounter),
    .io_input_toBuffer_0_ready(fetchBuffer_1_io_input_toBuffer_0_ready),
    .io_input_toBuffer_0_valid(fetchBuffer_1_io_input_toBuffer_0_valid),
    .io_input_toBuffer_0_bits_instruction(fetchBuffer_1_io_input_toBuffer_0_bits_instruction),
    .io_input_toBuffer_0_bits_programCounter(fetchBuffer_1_io_input_toBuffer_0_bits_programCounter),
    .io_input_empty(fetchBuffer_1_io_input_empty)
  );
  ReorderBuffer reorderBuffer_0 ( // @[B4Processor.scala 40:45]
    .clock(reorderBuffer_0_clock),
    .reset(reorderBuffer_0_reset),
    .io_decoders_0_source1_sourceRegister(reorderBuffer_0_io_decoders_0_source1_sourceRegister),
    .io_decoders_0_source1_matchingTag_valid(reorderBuffer_0_io_decoders_0_source1_matchingTag_valid),
    .io_decoders_0_source1_matchingTag_bits_id(reorderBuffer_0_io_decoders_0_source1_matchingTag_bits_id),
    .io_decoders_0_source1_value_valid(reorderBuffer_0_io_decoders_0_source1_value_valid),
    .io_decoders_0_source1_value_bits(reorderBuffer_0_io_decoders_0_source1_value_bits),
    .io_decoders_0_source2_sourceRegister(reorderBuffer_0_io_decoders_0_source2_sourceRegister),
    .io_decoders_0_source2_matchingTag_valid(reorderBuffer_0_io_decoders_0_source2_matchingTag_valid),
    .io_decoders_0_source2_matchingTag_bits_id(reorderBuffer_0_io_decoders_0_source2_matchingTag_bits_id),
    .io_decoders_0_source2_value_valid(reorderBuffer_0_io_decoders_0_source2_value_valid),
    .io_decoders_0_source2_value_bits(reorderBuffer_0_io_decoders_0_source2_value_bits),
    .io_decoders_0_destination_destinationRegister(reorderBuffer_0_io_decoders_0_destination_destinationRegister),
    .io_decoders_0_destination_destinationTag_id(reorderBuffer_0_io_decoders_0_destination_destinationTag_id),
    .io_decoders_0_destination_storeSign(reorderBuffer_0_io_decoders_0_destination_storeSign),
    .io_decoders_0_ready(reorderBuffer_0_io_decoders_0_ready),
    .io_decoders_0_valid(reorderBuffer_0_io_decoders_0_valid),
    .io_collectedOutputs_outputs_valid(reorderBuffer_0_io_collectedOutputs_outputs_valid),
    .io_collectedOutputs_outputs_bits_resultType(reorderBuffer_0_io_collectedOutputs_outputs_bits_resultType),
    .io_collectedOutputs_outputs_bits_value(reorderBuffer_0_io_collectedOutputs_outputs_bits_value),
    .io_collectedOutputs_outputs_bits_isError(reorderBuffer_0_io_collectedOutputs_outputs_bits_isError),
    .io_collectedOutputs_outputs_bits_tag_threadId(reorderBuffer_0_io_collectedOutputs_outputs_bits_tag_threadId),
    .io_collectedOutputs_outputs_bits_tag_id(reorderBuffer_0_io_collectedOutputs_outputs_bits_tag_id),
    .io_registerFile_0_valid(reorderBuffer_0_io_registerFile_0_valid),
    .io_registerFile_0_bits_destinationRegister(reorderBuffer_0_io_registerFile_0_bits_destinationRegister),
    .io_registerFile_0_bits_value(reorderBuffer_0_io_registerFile_0_bits_value),
    .io_registerFile_1_valid(reorderBuffer_0_io_registerFile_1_valid),
    .io_registerFile_1_bits_destinationRegister(reorderBuffer_0_io_registerFile_1_bits_destinationRegister),
    .io_registerFile_1_bits_value(reorderBuffer_0_io_registerFile_1_bits_value),
    .io_registerFile_2_valid(reorderBuffer_0_io_registerFile_2_valid),
    .io_registerFile_2_bits_destinationRegister(reorderBuffer_0_io_registerFile_2_bits_destinationRegister),
    .io_registerFile_2_bits_value(reorderBuffer_0_io_registerFile_2_bits_value),
    .io_registerFile_3_valid(reorderBuffer_0_io_registerFile_3_valid),
    .io_registerFile_3_bits_destinationRegister(reorderBuffer_0_io_registerFile_3_bits_destinationRegister),
    .io_registerFile_3_bits_value(reorderBuffer_0_io_registerFile_3_bits_value),
    .io_loadStoreQueue_0_valid(reorderBuffer_0_io_loadStoreQueue_0_valid),
    .io_loadStoreQueue_0_bits_destinationTag_id(reorderBuffer_0_io_loadStoreQueue_0_bits_destinationTag_id),
    .io_loadStoreQueue_1_valid(reorderBuffer_0_io_loadStoreQueue_1_valid),
    .io_loadStoreQueue_1_bits_destinationTag_id(reorderBuffer_0_io_loadStoreQueue_1_bits_destinationTag_id),
    .io_loadStoreQueue_2_valid(reorderBuffer_0_io_loadStoreQueue_2_valid),
    .io_loadStoreQueue_2_bits_destinationTag_id(reorderBuffer_0_io_loadStoreQueue_2_bits_destinationTag_id),
    .io_loadStoreQueue_3_valid(reorderBuffer_0_io_loadStoreQueue_3_valid),
    .io_loadStoreQueue_3_bits_destinationTag_id(reorderBuffer_0_io_loadStoreQueue_3_bits_destinationTag_id),
    .io_isEmpty(reorderBuffer_0_io_isEmpty),
    .io_csr_retireCount(reorderBuffer_0_io_csr_retireCount),
    .io_isError(reorderBuffer_0_io_isError)
  );
  ReorderBuffer_1 reorderBuffer_1 ( // @[B4Processor.scala 40:45]
    .clock(reorderBuffer_1_clock),
    .reset(reorderBuffer_1_reset),
    .io_decoders_0_source1_sourceRegister(reorderBuffer_1_io_decoders_0_source1_sourceRegister),
    .io_decoders_0_source1_matchingTag_valid(reorderBuffer_1_io_decoders_0_source1_matchingTag_valid),
    .io_decoders_0_source1_matchingTag_bits_id(reorderBuffer_1_io_decoders_0_source1_matchingTag_bits_id),
    .io_decoders_0_source1_value_valid(reorderBuffer_1_io_decoders_0_source1_value_valid),
    .io_decoders_0_source1_value_bits(reorderBuffer_1_io_decoders_0_source1_value_bits),
    .io_decoders_0_source2_sourceRegister(reorderBuffer_1_io_decoders_0_source2_sourceRegister),
    .io_decoders_0_source2_matchingTag_valid(reorderBuffer_1_io_decoders_0_source2_matchingTag_valid),
    .io_decoders_0_source2_matchingTag_bits_id(reorderBuffer_1_io_decoders_0_source2_matchingTag_bits_id),
    .io_decoders_0_source2_value_valid(reorderBuffer_1_io_decoders_0_source2_value_valid),
    .io_decoders_0_source2_value_bits(reorderBuffer_1_io_decoders_0_source2_value_bits),
    .io_decoders_0_destination_destinationRegister(reorderBuffer_1_io_decoders_0_destination_destinationRegister),
    .io_decoders_0_destination_destinationTag_id(reorderBuffer_1_io_decoders_0_destination_destinationTag_id),
    .io_decoders_0_destination_storeSign(reorderBuffer_1_io_decoders_0_destination_storeSign),
    .io_decoders_0_ready(reorderBuffer_1_io_decoders_0_ready),
    .io_decoders_0_valid(reorderBuffer_1_io_decoders_0_valid),
    .io_collectedOutputs_outputs_valid(reorderBuffer_1_io_collectedOutputs_outputs_valid),
    .io_collectedOutputs_outputs_bits_resultType(reorderBuffer_1_io_collectedOutputs_outputs_bits_resultType),
    .io_collectedOutputs_outputs_bits_value(reorderBuffer_1_io_collectedOutputs_outputs_bits_value),
    .io_collectedOutputs_outputs_bits_isError(reorderBuffer_1_io_collectedOutputs_outputs_bits_isError),
    .io_collectedOutputs_outputs_bits_tag_threadId(reorderBuffer_1_io_collectedOutputs_outputs_bits_tag_threadId),
    .io_collectedOutputs_outputs_bits_tag_id(reorderBuffer_1_io_collectedOutputs_outputs_bits_tag_id),
    .io_registerFile_0_valid(reorderBuffer_1_io_registerFile_0_valid),
    .io_registerFile_0_bits_destinationRegister(reorderBuffer_1_io_registerFile_0_bits_destinationRegister),
    .io_registerFile_0_bits_value(reorderBuffer_1_io_registerFile_0_bits_value),
    .io_registerFile_1_valid(reorderBuffer_1_io_registerFile_1_valid),
    .io_registerFile_1_bits_destinationRegister(reorderBuffer_1_io_registerFile_1_bits_destinationRegister),
    .io_registerFile_1_bits_value(reorderBuffer_1_io_registerFile_1_bits_value),
    .io_registerFile_2_valid(reorderBuffer_1_io_registerFile_2_valid),
    .io_registerFile_2_bits_destinationRegister(reorderBuffer_1_io_registerFile_2_bits_destinationRegister),
    .io_registerFile_2_bits_value(reorderBuffer_1_io_registerFile_2_bits_value),
    .io_registerFile_3_valid(reorderBuffer_1_io_registerFile_3_valid),
    .io_registerFile_3_bits_destinationRegister(reorderBuffer_1_io_registerFile_3_bits_destinationRegister),
    .io_registerFile_3_bits_value(reorderBuffer_1_io_registerFile_3_bits_value),
    .io_loadStoreQueue_0_valid(reorderBuffer_1_io_loadStoreQueue_0_valid),
    .io_loadStoreQueue_0_bits_destinationTag_id(reorderBuffer_1_io_loadStoreQueue_0_bits_destinationTag_id),
    .io_loadStoreQueue_1_valid(reorderBuffer_1_io_loadStoreQueue_1_valid),
    .io_loadStoreQueue_1_bits_destinationTag_id(reorderBuffer_1_io_loadStoreQueue_1_bits_destinationTag_id),
    .io_loadStoreQueue_2_valid(reorderBuffer_1_io_loadStoreQueue_2_valid),
    .io_loadStoreQueue_2_bits_destinationTag_id(reorderBuffer_1_io_loadStoreQueue_2_bits_destinationTag_id),
    .io_loadStoreQueue_3_valid(reorderBuffer_1_io_loadStoreQueue_3_valid),
    .io_loadStoreQueue_3_bits_destinationTag_id(reorderBuffer_1_io_loadStoreQueue_3_bits_destinationTag_id),
    .io_isEmpty(reorderBuffer_1_io_isEmpty),
    .io_csr_retireCount(reorderBuffer_1_io_csr_retireCount),
    .io_isError(reorderBuffer_1_io_isError)
  );
  RegisterFile registerFile_0 ( // @[B4Processor.scala 42:45]
    .clock(registerFile_0_clock),
    .reset(registerFile_0_reset),
    .io_decoders_0_sourceRegister1(registerFile_0_io_decoders_0_sourceRegister1),
    .io_decoders_0_sourceRegister2(registerFile_0_io_decoders_0_sourceRegister2),
    .io_decoders_0_value1(registerFile_0_io_decoders_0_value1),
    .io_decoders_0_value2(registerFile_0_io_decoders_0_value2),
    .io_reorderBuffer_0_valid(registerFile_0_io_reorderBuffer_0_valid),
    .io_reorderBuffer_0_bits_destinationRegister(registerFile_0_io_reorderBuffer_0_bits_destinationRegister),
    .io_reorderBuffer_0_bits_value(registerFile_0_io_reorderBuffer_0_bits_value),
    .io_reorderBuffer_1_valid(registerFile_0_io_reorderBuffer_1_valid),
    .io_reorderBuffer_1_bits_destinationRegister(registerFile_0_io_reorderBuffer_1_bits_destinationRegister),
    .io_reorderBuffer_1_bits_value(registerFile_0_io_reorderBuffer_1_bits_value),
    .io_reorderBuffer_2_valid(registerFile_0_io_reorderBuffer_2_valid),
    .io_reorderBuffer_2_bits_destinationRegister(registerFile_0_io_reorderBuffer_2_bits_destinationRegister),
    .io_reorderBuffer_2_bits_value(registerFile_0_io_reorderBuffer_2_bits_value),
    .io_reorderBuffer_3_valid(registerFile_0_io_reorderBuffer_3_valid),
    .io_reorderBuffer_3_bits_destinationRegister(registerFile_0_io_reorderBuffer_3_bits_destinationRegister),
    .io_reorderBuffer_3_bits_value(registerFile_0_io_reorderBuffer_3_bits_value)
  );
  RegisterFile_1 registerFile_1 ( // @[B4Processor.scala 42:45]
    .clock(registerFile_1_clock),
    .reset(registerFile_1_reset),
    .io_decoders_0_sourceRegister1(registerFile_1_io_decoders_0_sourceRegister1),
    .io_decoders_0_sourceRegister2(registerFile_1_io_decoders_0_sourceRegister2),
    .io_decoders_0_value1(registerFile_1_io_decoders_0_value1),
    .io_decoders_0_value2(registerFile_1_io_decoders_0_value2),
    .io_reorderBuffer_0_valid(registerFile_1_io_reorderBuffer_0_valid),
    .io_reorderBuffer_0_bits_destinationRegister(registerFile_1_io_reorderBuffer_0_bits_destinationRegister),
    .io_reorderBuffer_0_bits_value(registerFile_1_io_reorderBuffer_0_bits_value),
    .io_reorderBuffer_1_valid(registerFile_1_io_reorderBuffer_1_valid),
    .io_reorderBuffer_1_bits_destinationRegister(registerFile_1_io_reorderBuffer_1_bits_destinationRegister),
    .io_reorderBuffer_1_bits_value(registerFile_1_io_reorderBuffer_1_bits_value),
    .io_reorderBuffer_2_valid(registerFile_1_io_reorderBuffer_2_valid),
    .io_reorderBuffer_2_bits_destinationRegister(registerFile_1_io_reorderBuffer_2_bits_destinationRegister),
    .io_reorderBuffer_2_bits_value(registerFile_1_io_reorderBuffer_2_bits_value),
    .io_reorderBuffer_3_valid(registerFile_1_io_reorderBuffer_3_valid),
    .io_reorderBuffer_3_bits_destinationRegister(registerFile_1_io_reorderBuffer_3_bits_destinationRegister),
    .io_reorderBuffer_3_bits_value(registerFile_1_io_reorderBuffer_3_bits_value)
  );
  LoadStoreQueue loadStoreQueue_0 ( // @[B4Processor.scala 44:45]
    .clock(loadStoreQueue_0_clock),
    .reset(loadStoreQueue_0_reset),
    .io_decoders_0_ready(loadStoreQueue_0_io_decoders_0_ready),
    .io_decoders_0_valid(loadStoreQueue_0_io_decoders_0_valid),
    .io_decoders_0_bits_accessInfo_accessType(loadStoreQueue_0_io_decoders_0_bits_accessInfo_accessType),
    .io_decoders_0_bits_accessInfo_signed(loadStoreQueue_0_io_decoders_0_bits_accessInfo_signed),
    .io_decoders_0_bits_accessInfo_accessWidth(loadStoreQueue_0_io_decoders_0_bits_accessInfo_accessWidth),
    .io_decoders_0_bits_addressAndLoadResultTag_threadId(
      loadStoreQueue_0_io_decoders_0_bits_addressAndLoadResultTag_threadId),
    .io_decoders_0_bits_addressAndLoadResultTag_id(loadStoreQueue_0_io_decoders_0_bits_addressAndLoadResultTag_id),
    .io_decoders_0_bits_address(loadStoreQueue_0_io_decoders_0_bits_address),
    .io_decoders_0_bits_addressValid(loadStoreQueue_0_io_decoders_0_bits_addressValid),
    .io_decoders_0_bits_storeDataTag_threadId(loadStoreQueue_0_io_decoders_0_bits_storeDataTag_threadId),
    .io_decoders_0_bits_storeDataTag_id(loadStoreQueue_0_io_decoders_0_bits_storeDataTag_id),
    .io_decoders_0_bits_storeData(loadStoreQueue_0_io_decoders_0_bits_storeData),
    .io_decoders_0_bits_storeDataValid(loadStoreQueue_0_io_decoders_0_bits_storeDataValid),
    .io_outputCollector_outputs_valid(loadStoreQueue_0_io_outputCollector_outputs_valid),
    .io_outputCollector_outputs_bits_resultType(loadStoreQueue_0_io_outputCollector_outputs_bits_resultType),
    .io_outputCollector_outputs_bits_value(loadStoreQueue_0_io_outputCollector_outputs_bits_value),
    .io_outputCollector_outputs_bits_tag_threadId(loadStoreQueue_0_io_outputCollector_outputs_bits_tag_threadId),
    .io_outputCollector_outputs_bits_tag_id(loadStoreQueue_0_io_outputCollector_outputs_bits_tag_id),
    .io_reorderBuffer_0_valid(loadStoreQueue_0_io_reorderBuffer_0_valid),
    .io_reorderBuffer_0_bits_destinationTag_threadId(loadStoreQueue_0_io_reorderBuffer_0_bits_destinationTag_threadId),
    .io_reorderBuffer_0_bits_destinationTag_id(loadStoreQueue_0_io_reorderBuffer_0_bits_destinationTag_id),
    .io_reorderBuffer_1_valid(loadStoreQueue_0_io_reorderBuffer_1_valid),
    .io_reorderBuffer_1_bits_destinationTag_threadId(loadStoreQueue_0_io_reorderBuffer_1_bits_destinationTag_threadId),
    .io_reorderBuffer_1_bits_destinationTag_id(loadStoreQueue_0_io_reorderBuffer_1_bits_destinationTag_id),
    .io_reorderBuffer_2_valid(loadStoreQueue_0_io_reorderBuffer_2_valid),
    .io_reorderBuffer_2_bits_destinationTag_threadId(loadStoreQueue_0_io_reorderBuffer_2_bits_destinationTag_threadId),
    .io_reorderBuffer_2_bits_destinationTag_id(loadStoreQueue_0_io_reorderBuffer_2_bits_destinationTag_id),
    .io_reorderBuffer_3_valid(loadStoreQueue_0_io_reorderBuffer_3_valid),
    .io_reorderBuffer_3_bits_destinationTag_threadId(loadStoreQueue_0_io_reorderBuffer_3_bits_destinationTag_threadId),
    .io_reorderBuffer_3_bits_destinationTag_id(loadStoreQueue_0_io_reorderBuffer_3_bits_destinationTag_id),
    .io_memory_ready(loadStoreQueue_0_io_memory_ready),
    .io_memory_valid(loadStoreQueue_0_io_memory_valid),
    .io_memory_bits_address(loadStoreQueue_0_io_memory_bits_address),
    .io_memory_bits_tag_threadId(loadStoreQueue_0_io_memory_bits_tag_threadId),
    .io_memory_bits_tag_id(loadStoreQueue_0_io_memory_bits_tag_id),
    .io_memory_bits_data(loadStoreQueue_0_io_memory_bits_data),
    .io_memory_bits_accessInfo_accessType(loadStoreQueue_0_io_memory_bits_accessInfo_accessType),
    .io_memory_bits_accessInfo_signed(loadStoreQueue_0_io_memory_bits_accessInfo_signed),
    .io_memory_bits_accessInfo_accessWidth(loadStoreQueue_0_io_memory_bits_accessInfo_accessWidth),
    .io_isEmpty(loadStoreQueue_0_io_isEmpty)
  );
  LoadStoreQueue loadStoreQueue_1 ( // @[B4Processor.scala 44:45]
    .clock(loadStoreQueue_1_clock),
    .reset(loadStoreQueue_1_reset),
    .io_decoders_0_ready(loadStoreQueue_1_io_decoders_0_ready),
    .io_decoders_0_valid(loadStoreQueue_1_io_decoders_0_valid),
    .io_decoders_0_bits_accessInfo_accessType(loadStoreQueue_1_io_decoders_0_bits_accessInfo_accessType),
    .io_decoders_0_bits_accessInfo_signed(loadStoreQueue_1_io_decoders_0_bits_accessInfo_signed),
    .io_decoders_0_bits_accessInfo_accessWidth(loadStoreQueue_1_io_decoders_0_bits_accessInfo_accessWidth),
    .io_decoders_0_bits_addressAndLoadResultTag_threadId(
      loadStoreQueue_1_io_decoders_0_bits_addressAndLoadResultTag_threadId),
    .io_decoders_0_bits_addressAndLoadResultTag_id(loadStoreQueue_1_io_decoders_0_bits_addressAndLoadResultTag_id),
    .io_decoders_0_bits_address(loadStoreQueue_1_io_decoders_0_bits_address),
    .io_decoders_0_bits_addressValid(loadStoreQueue_1_io_decoders_0_bits_addressValid),
    .io_decoders_0_bits_storeDataTag_threadId(loadStoreQueue_1_io_decoders_0_bits_storeDataTag_threadId),
    .io_decoders_0_bits_storeDataTag_id(loadStoreQueue_1_io_decoders_0_bits_storeDataTag_id),
    .io_decoders_0_bits_storeData(loadStoreQueue_1_io_decoders_0_bits_storeData),
    .io_decoders_0_bits_storeDataValid(loadStoreQueue_1_io_decoders_0_bits_storeDataValid),
    .io_outputCollector_outputs_valid(loadStoreQueue_1_io_outputCollector_outputs_valid),
    .io_outputCollector_outputs_bits_resultType(loadStoreQueue_1_io_outputCollector_outputs_bits_resultType),
    .io_outputCollector_outputs_bits_value(loadStoreQueue_1_io_outputCollector_outputs_bits_value),
    .io_outputCollector_outputs_bits_tag_threadId(loadStoreQueue_1_io_outputCollector_outputs_bits_tag_threadId),
    .io_outputCollector_outputs_bits_tag_id(loadStoreQueue_1_io_outputCollector_outputs_bits_tag_id),
    .io_reorderBuffer_0_valid(loadStoreQueue_1_io_reorderBuffer_0_valid),
    .io_reorderBuffer_0_bits_destinationTag_threadId(loadStoreQueue_1_io_reorderBuffer_0_bits_destinationTag_threadId),
    .io_reorderBuffer_0_bits_destinationTag_id(loadStoreQueue_1_io_reorderBuffer_0_bits_destinationTag_id),
    .io_reorderBuffer_1_valid(loadStoreQueue_1_io_reorderBuffer_1_valid),
    .io_reorderBuffer_1_bits_destinationTag_threadId(loadStoreQueue_1_io_reorderBuffer_1_bits_destinationTag_threadId),
    .io_reorderBuffer_1_bits_destinationTag_id(loadStoreQueue_1_io_reorderBuffer_1_bits_destinationTag_id),
    .io_reorderBuffer_2_valid(loadStoreQueue_1_io_reorderBuffer_2_valid),
    .io_reorderBuffer_2_bits_destinationTag_threadId(loadStoreQueue_1_io_reorderBuffer_2_bits_destinationTag_threadId),
    .io_reorderBuffer_2_bits_destinationTag_id(loadStoreQueue_1_io_reorderBuffer_2_bits_destinationTag_id),
    .io_reorderBuffer_3_valid(loadStoreQueue_1_io_reorderBuffer_3_valid),
    .io_reorderBuffer_3_bits_destinationTag_threadId(loadStoreQueue_1_io_reorderBuffer_3_bits_destinationTag_threadId),
    .io_reorderBuffer_3_bits_destinationTag_id(loadStoreQueue_1_io_reorderBuffer_3_bits_destinationTag_id),
    .io_memory_ready(loadStoreQueue_1_io_memory_ready),
    .io_memory_valid(loadStoreQueue_1_io_memory_valid),
    .io_memory_bits_address(loadStoreQueue_1_io_memory_bits_address),
    .io_memory_bits_tag_threadId(loadStoreQueue_1_io_memory_bits_tag_threadId),
    .io_memory_bits_tag_id(loadStoreQueue_1_io_memory_bits_tag_id),
    .io_memory_bits_data(loadStoreQueue_1_io_memory_bits_data),
    .io_memory_bits_accessInfo_accessType(loadStoreQueue_1_io_memory_bits_accessInfo_accessType),
    .io_memory_bits_accessInfo_signed(loadStoreQueue_1_io_memory_bits_accessInfo_signed),
    .io_memory_bits_accessInfo_accessWidth(loadStoreQueue_1_io_memory_bits_accessInfo_accessWidth),
    .io_isEmpty(loadStoreQueue_1_io_isEmpty)
  );
  DataMemoryBuffer dataMemoryBuffer ( // @[B4Processor.scala 45:40]
    .clock(dataMemoryBuffer_clock),
    .reset(dataMemoryBuffer_reset),
    .io_dataIn_0_ready(dataMemoryBuffer_io_dataIn_0_ready),
    .io_dataIn_0_valid(dataMemoryBuffer_io_dataIn_0_valid),
    .io_dataIn_0_bits_address(dataMemoryBuffer_io_dataIn_0_bits_address),
    .io_dataIn_0_bits_tag_threadId(dataMemoryBuffer_io_dataIn_0_bits_tag_threadId),
    .io_dataIn_0_bits_tag_id(dataMemoryBuffer_io_dataIn_0_bits_tag_id),
    .io_dataIn_0_bits_data(dataMemoryBuffer_io_dataIn_0_bits_data),
    .io_dataIn_0_bits_accessInfo_accessType(dataMemoryBuffer_io_dataIn_0_bits_accessInfo_accessType),
    .io_dataIn_0_bits_accessInfo_signed(dataMemoryBuffer_io_dataIn_0_bits_accessInfo_signed),
    .io_dataIn_0_bits_accessInfo_accessWidth(dataMemoryBuffer_io_dataIn_0_bits_accessInfo_accessWidth),
    .io_dataIn_1_ready(dataMemoryBuffer_io_dataIn_1_ready),
    .io_dataIn_1_valid(dataMemoryBuffer_io_dataIn_1_valid),
    .io_dataIn_1_bits_address(dataMemoryBuffer_io_dataIn_1_bits_address),
    .io_dataIn_1_bits_tag_threadId(dataMemoryBuffer_io_dataIn_1_bits_tag_threadId),
    .io_dataIn_1_bits_tag_id(dataMemoryBuffer_io_dataIn_1_bits_tag_id),
    .io_dataIn_1_bits_data(dataMemoryBuffer_io_dataIn_1_bits_data),
    .io_dataIn_1_bits_accessInfo_accessType(dataMemoryBuffer_io_dataIn_1_bits_accessInfo_accessType),
    .io_dataIn_1_bits_accessInfo_signed(dataMemoryBuffer_io_dataIn_1_bits_accessInfo_signed),
    .io_dataIn_1_bits_accessInfo_accessWidth(dataMemoryBuffer_io_dataIn_1_bits_accessInfo_accessWidth),
    .io_dataReadRequest_ready(dataMemoryBuffer_io_dataReadRequest_ready),
    .io_dataReadRequest_valid(dataMemoryBuffer_io_dataReadRequest_valid),
    .io_dataReadRequest_bits_address(dataMemoryBuffer_io_dataReadRequest_bits_address),
    .io_dataReadRequest_bits_size(dataMemoryBuffer_io_dataReadRequest_bits_size),
    .io_dataReadRequest_bits_signed(dataMemoryBuffer_io_dataReadRequest_bits_signed),
    .io_dataReadRequest_bits_outputTag_threadId(dataMemoryBuffer_io_dataReadRequest_bits_outputTag_threadId),
    .io_dataReadRequest_bits_outputTag_id(dataMemoryBuffer_io_dataReadRequest_bits_outputTag_id),
    .io_dataWriteRequest_ready(dataMemoryBuffer_io_dataWriteRequest_ready),
    .io_dataWriteRequest_valid(dataMemoryBuffer_io_dataWriteRequest_valid),
    .io_dataWriteRequest_bits_address(dataMemoryBuffer_io_dataWriteRequest_bits_address),
    .io_dataWriteRequest_bits_data(dataMemoryBuffer_io_dataWriteRequest_bits_data),
    .io_dataWriteRequest_bits_mask(dataMemoryBuffer_io_dataWriteRequest_bits_mask)
  );
  OutputCollector outputCollector ( // @[B4Processor.scala 47:31]
    .clock(outputCollector_clock),
    .reset(outputCollector_reset),
    .io_outputs_0_outputs_valid(outputCollector_io_outputs_0_outputs_valid),
    .io_outputs_0_outputs_bits_resultType(outputCollector_io_outputs_0_outputs_bits_resultType),
    .io_outputs_0_outputs_bits_value(outputCollector_io_outputs_0_outputs_bits_value),
    .io_outputs_0_outputs_bits_isError(outputCollector_io_outputs_0_outputs_bits_isError),
    .io_outputs_0_outputs_bits_tag_threadId(outputCollector_io_outputs_0_outputs_bits_tag_threadId),
    .io_outputs_0_outputs_bits_tag_id(outputCollector_io_outputs_0_outputs_bits_tag_id),
    .io_outputs_1_outputs_valid(outputCollector_io_outputs_1_outputs_valid),
    .io_outputs_1_outputs_bits_resultType(outputCollector_io_outputs_1_outputs_bits_resultType),
    .io_outputs_1_outputs_bits_value(outputCollector_io_outputs_1_outputs_bits_value),
    .io_outputs_1_outputs_bits_isError(outputCollector_io_outputs_1_outputs_bits_isError),
    .io_outputs_1_outputs_bits_tag_threadId(outputCollector_io_outputs_1_outputs_bits_tag_threadId),
    .io_outputs_1_outputs_bits_tag_id(outputCollector_io_outputs_1_outputs_bits_tag_id),
    .io_executor_0_ready(outputCollector_io_executor_0_ready),
    .io_executor_0_valid(outputCollector_io_executor_0_valid),
    .io_executor_0_bits_resultType(outputCollector_io_executor_0_bits_resultType),
    .io_executor_0_bits_value(outputCollector_io_executor_0_bits_value),
    .io_executor_0_bits_tag_threadId(outputCollector_io_executor_0_bits_tag_threadId),
    .io_executor_0_bits_tag_id(outputCollector_io_executor_0_bits_tag_id),
    .io_executor_1_ready(outputCollector_io_executor_1_ready),
    .io_executor_1_valid(outputCollector_io_executor_1_valid),
    .io_executor_1_bits_resultType(outputCollector_io_executor_1_bits_resultType),
    .io_executor_1_bits_value(outputCollector_io_executor_1_bits_value),
    .io_executor_1_bits_tag_threadId(outputCollector_io_executor_1_bits_tag_threadId),
    .io_executor_1_bits_tag_id(outputCollector_io_executor_1_bits_tag_id),
    .io_dataMemory_ready(outputCollector_io_dataMemory_ready),
    .io_dataMemory_valid(outputCollector_io_dataMemory_valid),
    .io_dataMemory_bits_value(outputCollector_io_dataMemory_bits_value),
    .io_dataMemory_bits_isError(outputCollector_io_dataMemory_bits_isError),
    .io_dataMemory_bits_tag_threadId(outputCollector_io_dataMemory_bits_tag_threadId),
    .io_dataMemory_bits_tag_id(outputCollector_io_dataMemory_bits_tag_id),
    .io_csr_0_ready(outputCollector_io_csr_0_ready),
    .io_csr_0_valid(outputCollector_io_csr_0_valid),
    .io_csr_0_bits_value(outputCollector_io_csr_0_bits_value),
    .io_csr_0_bits_isError(outputCollector_io_csr_0_bits_isError),
    .io_csr_0_bits_tag_threadId(outputCollector_io_csr_0_bits_tag_threadId),
    .io_csr_0_bits_tag_id(outputCollector_io_csr_0_bits_tag_id),
    .io_csr_1_ready(outputCollector_io_csr_1_ready),
    .io_csr_1_valid(outputCollector_io_csr_1_valid),
    .io_csr_1_bits_value(outputCollector_io_csr_1_bits_value),
    .io_csr_1_bits_isError(outputCollector_io_csr_1_bits_isError),
    .io_csr_1_bits_tag_threadId(outputCollector_io_csr_1_bits_tag_threadId),
    .io_csr_1_bits_tag_id(outputCollector_io_csr_1_bits_tag_id),
    .io_isError_0(outputCollector_io_isError_0),
    .io_isError_1(outputCollector_io_isError_1)
  );
  BranchOutputCollector branchAddressCollector ( // @[B4Processor.scala 48:46]
    .clock(branchAddressCollector_clock),
    .reset(branchAddressCollector_reset),
    .io_fetch_0_addresses_valid(branchAddressCollector_io_fetch_0_addresses_valid),
    .io_fetch_0_addresses_bits_threadId(branchAddressCollector_io_fetch_0_addresses_bits_threadId),
    .io_fetch_0_addresses_bits_programCounterOffset(
      branchAddressCollector_io_fetch_0_addresses_bits_programCounterOffset),
    .io_fetch_1_addresses_valid(branchAddressCollector_io_fetch_1_addresses_valid),
    .io_fetch_1_addresses_bits_threadId(branchAddressCollector_io_fetch_1_addresses_bits_threadId),
    .io_fetch_1_addresses_bits_programCounterOffset(
      branchAddressCollector_io_fetch_1_addresses_bits_programCounterOffset),
    .io_executor_0_ready(branchAddressCollector_io_executor_0_ready),
    .io_executor_0_valid(branchAddressCollector_io_executor_0_valid),
    .io_executor_0_bits_threadId(branchAddressCollector_io_executor_0_bits_threadId),
    .io_executor_0_bits_programCounterOffset(branchAddressCollector_io_executor_0_bits_programCounterOffset),
    .io_executor_1_ready(branchAddressCollector_io_executor_1_ready),
    .io_executor_1_valid(branchAddressCollector_io_executor_1_valid),
    .io_executor_1_bits_threadId(branchAddressCollector_io_executor_1_bits_threadId),
    .io_executor_1_bits_programCounterOffset(branchAddressCollector_io_executor_1_bits_programCounterOffset),
    .io_isError_0(branchAddressCollector_io_isError_0),
    .io_isError_1(branchAddressCollector_io_isError_1)
  );
  Uncompresser uncompresser_0_0 ( // @[B4Processor.scala 51:45]
    .io_fetch_ready(uncompresser_0_0_io_fetch_ready),
    .io_fetch_valid(uncompresser_0_0_io_fetch_valid),
    .io_fetch_bits_instruction(uncompresser_0_0_io_fetch_bits_instruction),
    .io_fetch_bits_programCounter(uncompresser_0_0_io_fetch_bits_programCounter),
    .io_decoder_ready(uncompresser_0_0_io_decoder_ready),
    .io_decoder_valid(uncompresser_0_0_io_decoder_valid),
    .io_decoder_bits_instruction(uncompresser_0_0_io_decoder_bits_instruction),
    .io_decoder_bits_programCounter(uncompresser_0_0_io_decoder_bits_programCounter),
    .io_decoder_bits_wasCompressed(uncompresser_0_0_io_decoder_bits_wasCompressed)
  );
  Uncompresser uncompresser_1_0 ( // @[B4Processor.scala 51:45]
    .io_fetch_ready(uncompresser_1_0_io_fetch_ready),
    .io_fetch_valid(uncompresser_1_0_io_fetch_valid),
    .io_fetch_bits_instruction(uncompresser_1_0_io_fetch_bits_instruction),
    .io_fetch_bits_programCounter(uncompresser_1_0_io_fetch_bits_programCounter),
    .io_decoder_ready(uncompresser_1_0_io_decoder_ready),
    .io_decoder_valid(uncompresser_1_0_io_decoder_valid),
    .io_decoder_bits_instruction(uncompresser_1_0_io_decoder_bits_instruction),
    .io_decoder_bits_programCounter(uncompresser_1_0_io_decoder_bits_programCounter),
    .io_decoder_bits_wasCompressed(uncompresser_1_0_io_decoder_bits_wasCompressed)
  );
  Decoder decoders_0_0 ( // @[B4Processor.scala 54:54]
    .io_instructionFetch_ready(decoders_0_0_io_instructionFetch_ready),
    .io_instructionFetch_valid(decoders_0_0_io_instructionFetch_valid),
    .io_instructionFetch_bits_instruction(decoders_0_0_io_instructionFetch_bits_instruction),
    .io_instructionFetch_bits_programCounter(decoders_0_0_io_instructionFetch_bits_programCounter),
    .io_instructionFetch_bits_wasCompressed(decoders_0_0_io_instructionFetch_bits_wasCompressed),
    .io_reorderBuffer_source1_sourceRegister(decoders_0_0_io_reorderBuffer_source1_sourceRegister),
    .io_reorderBuffer_source1_matchingTag_valid(decoders_0_0_io_reorderBuffer_source1_matchingTag_valid),
    .io_reorderBuffer_source1_matchingTag_bits_id(decoders_0_0_io_reorderBuffer_source1_matchingTag_bits_id),
    .io_reorderBuffer_source1_value_valid(decoders_0_0_io_reorderBuffer_source1_value_valid),
    .io_reorderBuffer_source1_value_bits(decoders_0_0_io_reorderBuffer_source1_value_bits),
    .io_reorderBuffer_source2_sourceRegister(decoders_0_0_io_reorderBuffer_source2_sourceRegister),
    .io_reorderBuffer_source2_matchingTag_valid(decoders_0_0_io_reorderBuffer_source2_matchingTag_valid),
    .io_reorderBuffer_source2_matchingTag_bits_id(decoders_0_0_io_reorderBuffer_source2_matchingTag_bits_id),
    .io_reorderBuffer_source2_value_valid(decoders_0_0_io_reorderBuffer_source2_value_valid),
    .io_reorderBuffer_source2_value_bits(decoders_0_0_io_reorderBuffer_source2_value_bits),
    .io_reorderBuffer_destination_destinationRegister(decoders_0_0_io_reorderBuffer_destination_destinationRegister),
    .io_reorderBuffer_destination_destinationTag_id(decoders_0_0_io_reorderBuffer_destination_destinationTag_id),
    .io_reorderBuffer_destination_storeSign(decoders_0_0_io_reorderBuffer_destination_storeSign),
    .io_reorderBuffer_ready(decoders_0_0_io_reorderBuffer_ready),
    .io_reorderBuffer_valid(decoders_0_0_io_reorderBuffer_valid),
    .io_outputCollector_outputs_valid(decoders_0_0_io_outputCollector_outputs_valid),
    .io_outputCollector_outputs_bits_resultType(decoders_0_0_io_outputCollector_outputs_bits_resultType),
    .io_outputCollector_outputs_bits_value(decoders_0_0_io_outputCollector_outputs_bits_value),
    .io_outputCollector_outputs_bits_tag_threadId(decoders_0_0_io_outputCollector_outputs_bits_tag_threadId),
    .io_outputCollector_outputs_bits_tag_id(decoders_0_0_io_outputCollector_outputs_bits_tag_id),
    .io_registerFile_sourceRegister1(decoders_0_0_io_registerFile_sourceRegister1),
    .io_registerFile_sourceRegister2(decoders_0_0_io_registerFile_sourceRegister2),
    .io_registerFile_value1(decoders_0_0_io_registerFile_value1),
    .io_registerFile_value2(decoders_0_0_io_registerFile_value2),
    .io_reservationStation_ready(decoders_0_0_io_reservationStation_ready),
    .io_reservationStation_entry_opcode(decoders_0_0_io_reservationStation_entry_opcode),
    .io_reservationStation_entry_function3(decoders_0_0_io_reservationStation_entry_function3),
    .io_reservationStation_entry_immediateOrFunction7(decoders_0_0_io_reservationStation_entry_immediateOrFunction7),
    .io_reservationStation_entry_sourceTag1_threadId(decoders_0_0_io_reservationStation_entry_sourceTag1_threadId),
    .io_reservationStation_entry_sourceTag1_id(decoders_0_0_io_reservationStation_entry_sourceTag1_id),
    .io_reservationStation_entry_ready1(decoders_0_0_io_reservationStation_entry_ready1),
    .io_reservationStation_entry_value1(decoders_0_0_io_reservationStation_entry_value1),
    .io_reservationStation_entry_sourceTag2_threadId(decoders_0_0_io_reservationStation_entry_sourceTag2_threadId),
    .io_reservationStation_entry_sourceTag2_id(decoders_0_0_io_reservationStation_entry_sourceTag2_id),
    .io_reservationStation_entry_ready2(decoders_0_0_io_reservationStation_entry_ready2),
    .io_reservationStation_entry_value2(decoders_0_0_io_reservationStation_entry_value2),
    .io_reservationStation_entry_destinationTag_threadId(
      decoders_0_0_io_reservationStation_entry_destinationTag_threadId),
    .io_reservationStation_entry_destinationTag_id(decoders_0_0_io_reservationStation_entry_destinationTag_id),
    .io_reservationStation_entry_wasCompressed(decoders_0_0_io_reservationStation_entry_wasCompressed),
    .io_reservationStation_entry_valid(decoders_0_0_io_reservationStation_entry_valid),
    .io_loadStoreQueue_ready(decoders_0_0_io_loadStoreQueue_ready),
    .io_loadStoreQueue_valid(decoders_0_0_io_loadStoreQueue_valid),
    .io_loadStoreQueue_bits_accessInfo_accessType(decoders_0_0_io_loadStoreQueue_bits_accessInfo_accessType),
    .io_loadStoreQueue_bits_accessInfo_signed(decoders_0_0_io_loadStoreQueue_bits_accessInfo_signed),
    .io_loadStoreQueue_bits_accessInfo_accessWidth(decoders_0_0_io_loadStoreQueue_bits_accessInfo_accessWidth),
    .io_loadStoreQueue_bits_addressAndLoadResultTag_threadId(
      decoders_0_0_io_loadStoreQueue_bits_addressAndLoadResultTag_threadId),
    .io_loadStoreQueue_bits_addressAndLoadResultTag_id(decoders_0_0_io_loadStoreQueue_bits_addressAndLoadResultTag_id),
    .io_loadStoreQueue_bits_address(decoders_0_0_io_loadStoreQueue_bits_address),
    .io_loadStoreQueue_bits_addressValid(decoders_0_0_io_loadStoreQueue_bits_addressValid),
    .io_loadStoreQueue_bits_storeDataTag_threadId(decoders_0_0_io_loadStoreQueue_bits_storeDataTag_threadId),
    .io_loadStoreQueue_bits_storeDataTag_id(decoders_0_0_io_loadStoreQueue_bits_storeDataTag_id),
    .io_loadStoreQueue_bits_storeData(decoders_0_0_io_loadStoreQueue_bits_storeData),
    .io_loadStoreQueue_bits_storeDataValid(decoders_0_0_io_loadStoreQueue_bits_storeDataValid),
    .io_csr_ready(decoders_0_0_io_csr_ready),
    .io_csr_valid(decoders_0_0_io_csr_valid),
    .io_csr_bits_sourceTag_threadId(decoders_0_0_io_csr_bits_sourceTag_threadId),
    .io_csr_bits_sourceTag_id(decoders_0_0_io_csr_bits_sourceTag_id),
    .io_csr_bits_destinationTag_id(decoders_0_0_io_csr_bits_destinationTag_id),
    .io_csr_bits_value(decoders_0_0_io_csr_bits_value),
    .io_csr_bits_ready(decoders_0_0_io_csr_bits_ready),
    .io_csr_bits_address(decoders_0_0_io_csr_bits_address),
    .io_csr_bits_csrAccessType(decoders_0_0_io_csr_bits_csrAccessType)
  );
  Decoder_1 decoders_1_0 ( // @[B4Processor.scala 54:54]
    .io_instructionFetch_ready(decoders_1_0_io_instructionFetch_ready),
    .io_instructionFetch_valid(decoders_1_0_io_instructionFetch_valid),
    .io_instructionFetch_bits_instruction(decoders_1_0_io_instructionFetch_bits_instruction),
    .io_instructionFetch_bits_programCounter(decoders_1_0_io_instructionFetch_bits_programCounter),
    .io_instructionFetch_bits_wasCompressed(decoders_1_0_io_instructionFetch_bits_wasCompressed),
    .io_reorderBuffer_source1_sourceRegister(decoders_1_0_io_reorderBuffer_source1_sourceRegister),
    .io_reorderBuffer_source1_matchingTag_valid(decoders_1_0_io_reorderBuffer_source1_matchingTag_valid),
    .io_reorderBuffer_source1_matchingTag_bits_id(decoders_1_0_io_reorderBuffer_source1_matchingTag_bits_id),
    .io_reorderBuffer_source1_value_valid(decoders_1_0_io_reorderBuffer_source1_value_valid),
    .io_reorderBuffer_source1_value_bits(decoders_1_0_io_reorderBuffer_source1_value_bits),
    .io_reorderBuffer_source2_sourceRegister(decoders_1_0_io_reorderBuffer_source2_sourceRegister),
    .io_reorderBuffer_source2_matchingTag_valid(decoders_1_0_io_reorderBuffer_source2_matchingTag_valid),
    .io_reorderBuffer_source2_matchingTag_bits_id(decoders_1_0_io_reorderBuffer_source2_matchingTag_bits_id),
    .io_reorderBuffer_source2_value_valid(decoders_1_0_io_reorderBuffer_source2_value_valid),
    .io_reorderBuffer_source2_value_bits(decoders_1_0_io_reorderBuffer_source2_value_bits),
    .io_reorderBuffer_destination_destinationRegister(decoders_1_0_io_reorderBuffer_destination_destinationRegister),
    .io_reorderBuffer_destination_destinationTag_id(decoders_1_0_io_reorderBuffer_destination_destinationTag_id),
    .io_reorderBuffer_destination_storeSign(decoders_1_0_io_reorderBuffer_destination_storeSign),
    .io_reorderBuffer_ready(decoders_1_0_io_reorderBuffer_ready),
    .io_reorderBuffer_valid(decoders_1_0_io_reorderBuffer_valid),
    .io_outputCollector_outputs_valid(decoders_1_0_io_outputCollector_outputs_valid),
    .io_outputCollector_outputs_bits_resultType(decoders_1_0_io_outputCollector_outputs_bits_resultType),
    .io_outputCollector_outputs_bits_value(decoders_1_0_io_outputCollector_outputs_bits_value),
    .io_outputCollector_outputs_bits_tag_threadId(decoders_1_0_io_outputCollector_outputs_bits_tag_threadId),
    .io_outputCollector_outputs_bits_tag_id(decoders_1_0_io_outputCollector_outputs_bits_tag_id),
    .io_registerFile_sourceRegister1(decoders_1_0_io_registerFile_sourceRegister1),
    .io_registerFile_sourceRegister2(decoders_1_0_io_registerFile_sourceRegister2),
    .io_registerFile_value1(decoders_1_0_io_registerFile_value1),
    .io_registerFile_value2(decoders_1_0_io_registerFile_value2),
    .io_reservationStation_ready(decoders_1_0_io_reservationStation_ready),
    .io_reservationStation_entry_opcode(decoders_1_0_io_reservationStation_entry_opcode),
    .io_reservationStation_entry_function3(decoders_1_0_io_reservationStation_entry_function3),
    .io_reservationStation_entry_immediateOrFunction7(decoders_1_0_io_reservationStation_entry_immediateOrFunction7),
    .io_reservationStation_entry_sourceTag1_threadId(decoders_1_0_io_reservationStation_entry_sourceTag1_threadId),
    .io_reservationStation_entry_sourceTag1_id(decoders_1_0_io_reservationStation_entry_sourceTag1_id),
    .io_reservationStation_entry_ready1(decoders_1_0_io_reservationStation_entry_ready1),
    .io_reservationStation_entry_value1(decoders_1_0_io_reservationStation_entry_value1),
    .io_reservationStation_entry_sourceTag2_threadId(decoders_1_0_io_reservationStation_entry_sourceTag2_threadId),
    .io_reservationStation_entry_sourceTag2_id(decoders_1_0_io_reservationStation_entry_sourceTag2_id),
    .io_reservationStation_entry_ready2(decoders_1_0_io_reservationStation_entry_ready2),
    .io_reservationStation_entry_value2(decoders_1_0_io_reservationStation_entry_value2),
    .io_reservationStation_entry_destinationTag_threadId(
      decoders_1_0_io_reservationStation_entry_destinationTag_threadId),
    .io_reservationStation_entry_destinationTag_id(decoders_1_0_io_reservationStation_entry_destinationTag_id),
    .io_reservationStation_entry_wasCompressed(decoders_1_0_io_reservationStation_entry_wasCompressed),
    .io_reservationStation_entry_valid(decoders_1_0_io_reservationStation_entry_valid),
    .io_loadStoreQueue_ready(decoders_1_0_io_loadStoreQueue_ready),
    .io_loadStoreQueue_valid(decoders_1_0_io_loadStoreQueue_valid),
    .io_loadStoreQueue_bits_accessInfo_accessType(decoders_1_0_io_loadStoreQueue_bits_accessInfo_accessType),
    .io_loadStoreQueue_bits_accessInfo_signed(decoders_1_0_io_loadStoreQueue_bits_accessInfo_signed),
    .io_loadStoreQueue_bits_accessInfo_accessWidth(decoders_1_0_io_loadStoreQueue_bits_accessInfo_accessWidth),
    .io_loadStoreQueue_bits_addressAndLoadResultTag_threadId(
      decoders_1_0_io_loadStoreQueue_bits_addressAndLoadResultTag_threadId),
    .io_loadStoreQueue_bits_addressAndLoadResultTag_id(decoders_1_0_io_loadStoreQueue_bits_addressAndLoadResultTag_id),
    .io_loadStoreQueue_bits_address(decoders_1_0_io_loadStoreQueue_bits_address),
    .io_loadStoreQueue_bits_addressValid(decoders_1_0_io_loadStoreQueue_bits_addressValid),
    .io_loadStoreQueue_bits_storeDataTag_threadId(decoders_1_0_io_loadStoreQueue_bits_storeDataTag_threadId),
    .io_loadStoreQueue_bits_storeDataTag_id(decoders_1_0_io_loadStoreQueue_bits_storeDataTag_id),
    .io_loadStoreQueue_bits_storeData(decoders_1_0_io_loadStoreQueue_bits_storeData),
    .io_loadStoreQueue_bits_storeDataValid(decoders_1_0_io_loadStoreQueue_bits_storeDataValid),
    .io_csr_ready(decoders_1_0_io_csr_ready),
    .io_csr_valid(decoders_1_0_io_csr_valid),
    .io_csr_bits_sourceTag_threadId(decoders_1_0_io_csr_bits_sourceTag_threadId),
    .io_csr_bits_sourceTag_id(decoders_1_0_io_csr_bits_sourceTag_id),
    .io_csr_bits_destinationTag_id(decoders_1_0_io_csr_bits_destinationTag_id),
    .io_csr_bits_value(decoders_1_0_io_csr_bits_value),
    .io_csr_bits_ready(decoders_1_0_io_csr_bits_ready),
    .io_csr_bits_address(decoders_1_0_io_csr_bits_address),
    .io_csr_bits_csrAccessType(decoders_1_0_io_csr_bits_csrAccessType)
  );
  ReservationStation reservationStation ( // @[B4Processor.scala 56:42]
    .clock(reservationStation_clock),
    .reset(reservationStation_reset),
    .io_collectedOutput_0_outputs_valid(reservationStation_io_collectedOutput_0_outputs_valid),
    .io_collectedOutput_0_outputs_bits_resultType(reservationStation_io_collectedOutput_0_outputs_bits_resultType),
    .io_collectedOutput_0_outputs_bits_value(reservationStation_io_collectedOutput_0_outputs_bits_value),
    .io_collectedOutput_0_outputs_bits_tag_threadId(reservationStation_io_collectedOutput_0_outputs_bits_tag_threadId),
    .io_collectedOutput_0_outputs_bits_tag_id(reservationStation_io_collectedOutput_0_outputs_bits_tag_id),
    .io_collectedOutput_1_outputs_valid(reservationStation_io_collectedOutput_1_outputs_valid),
    .io_collectedOutput_1_outputs_bits_resultType(reservationStation_io_collectedOutput_1_outputs_bits_resultType),
    .io_collectedOutput_1_outputs_bits_value(reservationStation_io_collectedOutput_1_outputs_bits_value),
    .io_collectedOutput_1_outputs_bits_tag_threadId(reservationStation_io_collectedOutput_1_outputs_bits_tag_threadId),
    .io_collectedOutput_1_outputs_bits_tag_id(reservationStation_io_collectedOutput_1_outputs_bits_tag_id),
    .io_executor_0_ready(reservationStation_io_executor_0_ready),
    .io_executor_0_valid(reservationStation_io_executor_0_valid),
    .io_executor_0_bits_destinationTag_threadId(reservationStation_io_executor_0_bits_destinationTag_threadId),
    .io_executor_0_bits_destinationTag_id(reservationStation_io_executor_0_bits_destinationTag_id),
    .io_executor_0_bits_value1(reservationStation_io_executor_0_bits_value1),
    .io_executor_0_bits_value2(reservationStation_io_executor_0_bits_value2),
    .io_executor_0_bits_function3(reservationStation_io_executor_0_bits_function3),
    .io_executor_0_bits_immediateOrFunction7(reservationStation_io_executor_0_bits_immediateOrFunction7),
    .io_executor_0_bits_opcode(reservationStation_io_executor_0_bits_opcode),
    .io_executor_0_bits_wasCompressed(reservationStation_io_executor_0_bits_wasCompressed),
    .io_executor_1_ready(reservationStation_io_executor_1_ready),
    .io_executor_1_valid(reservationStation_io_executor_1_valid),
    .io_executor_1_bits_destinationTag_threadId(reservationStation_io_executor_1_bits_destinationTag_threadId),
    .io_executor_1_bits_destinationTag_id(reservationStation_io_executor_1_bits_destinationTag_id),
    .io_executor_1_bits_value1(reservationStation_io_executor_1_bits_value1),
    .io_executor_1_bits_value2(reservationStation_io_executor_1_bits_value2),
    .io_executor_1_bits_function3(reservationStation_io_executor_1_bits_function3),
    .io_executor_1_bits_immediateOrFunction7(reservationStation_io_executor_1_bits_immediateOrFunction7),
    .io_executor_1_bits_opcode(reservationStation_io_executor_1_bits_opcode),
    .io_executor_1_bits_wasCompressed(reservationStation_io_executor_1_bits_wasCompressed),
    .io_decoder_0_ready(reservationStation_io_decoder_0_ready),
    .io_decoder_0_entry_opcode(reservationStation_io_decoder_0_entry_opcode),
    .io_decoder_0_entry_function3(reservationStation_io_decoder_0_entry_function3),
    .io_decoder_0_entry_immediateOrFunction7(reservationStation_io_decoder_0_entry_immediateOrFunction7),
    .io_decoder_0_entry_sourceTag1_threadId(reservationStation_io_decoder_0_entry_sourceTag1_threadId),
    .io_decoder_0_entry_sourceTag1_id(reservationStation_io_decoder_0_entry_sourceTag1_id),
    .io_decoder_0_entry_ready1(reservationStation_io_decoder_0_entry_ready1),
    .io_decoder_0_entry_value1(reservationStation_io_decoder_0_entry_value1),
    .io_decoder_0_entry_sourceTag2_threadId(reservationStation_io_decoder_0_entry_sourceTag2_threadId),
    .io_decoder_0_entry_sourceTag2_id(reservationStation_io_decoder_0_entry_sourceTag2_id),
    .io_decoder_0_entry_ready2(reservationStation_io_decoder_0_entry_ready2),
    .io_decoder_0_entry_value2(reservationStation_io_decoder_0_entry_value2),
    .io_decoder_0_entry_destinationTag_id(reservationStation_io_decoder_0_entry_destinationTag_id),
    .io_decoder_0_entry_wasCompressed(reservationStation_io_decoder_0_entry_wasCompressed),
    .io_decoder_0_entry_valid(reservationStation_io_decoder_0_entry_valid),
    .io_decoder_1_ready(reservationStation_io_decoder_1_ready),
    .io_decoder_1_entry_opcode(reservationStation_io_decoder_1_entry_opcode),
    .io_decoder_1_entry_function3(reservationStation_io_decoder_1_entry_function3),
    .io_decoder_1_entry_immediateOrFunction7(reservationStation_io_decoder_1_entry_immediateOrFunction7),
    .io_decoder_1_entry_sourceTag1_threadId(reservationStation_io_decoder_1_entry_sourceTag1_threadId),
    .io_decoder_1_entry_sourceTag1_id(reservationStation_io_decoder_1_entry_sourceTag1_id),
    .io_decoder_1_entry_ready1(reservationStation_io_decoder_1_entry_ready1),
    .io_decoder_1_entry_value1(reservationStation_io_decoder_1_entry_value1),
    .io_decoder_1_entry_sourceTag2_threadId(reservationStation_io_decoder_1_entry_sourceTag2_threadId),
    .io_decoder_1_entry_sourceTag2_id(reservationStation_io_decoder_1_entry_sourceTag2_id),
    .io_decoder_1_entry_ready2(reservationStation_io_decoder_1_entry_ready2),
    .io_decoder_1_entry_value2(reservationStation_io_decoder_1_entry_value2),
    .io_decoder_1_entry_destinationTag_id(reservationStation_io_decoder_1_entry_destinationTag_id),
    .io_decoder_1_entry_wasCompressed(reservationStation_io_decoder_1_entry_wasCompressed),
    .io_decoder_1_entry_valid(reservationStation_io_decoder_1_entry_valid)
  );
  Executor executors_0 ( // @[B4Processor.scala 57:60]
    .io_reservationStation_ready(executors_0_io_reservationStation_ready),
    .io_reservationStation_valid(executors_0_io_reservationStation_valid),
    .io_reservationStation_bits_destinationTag_threadId(executors_0_io_reservationStation_bits_destinationTag_threadId),
    .io_reservationStation_bits_destinationTag_id(executors_0_io_reservationStation_bits_destinationTag_id),
    .io_reservationStation_bits_value1(executors_0_io_reservationStation_bits_value1),
    .io_reservationStation_bits_value2(executors_0_io_reservationStation_bits_value2),
    .io_reservationStation_bits_function3(executors_0_io_reservationStation_bits_function3),
    .io_reservationStation_bits_immediateOrFunction7(executors_0_io_reservationStation_bits_immediateOrFunction7),
    .io_reservationStation_bits_opcode(executors_0_io_reservationStation_bits_opcode),
    .io_reservationStation_bits_wasCompressed(executors_0_io_reservationStation_bits_wasCompressed),
    .io_out_ready(executors_0_io_out_ready),
    .io_out_valid(executors_0_io_out_valid),
    .io_out_bits_resultType(executors_0_io_out_bits_resultType),
    .io_out_bits_value(executors_0_io_out_bits_value),
    .io_out_bits_tag_threadId(executors_0_io_out_bits_tag_threadId),
    .io_out_bits_tag_id(executors_0_io_out_bits_tag_id),
    .io_fetch_ready(executors_0_io_fetch_ready),
    .io_fetch_valid(executors_0_io_fetch_valid),
    .io_fetch_bits_threadId(executors_0_io_fetch_bits_threadId),
    .io_fetch_bits_programCounterOffset(executors_0_io_fetch_bits_programCounterOffset)
  );
  Executor executors_1 ( // @[B4Processor.scala 57:60]
    .io_reservationStation_ready(executors_1_io_reservationStation_ready),
    .io_reservationStation_valid(executors_1_io_reservationStation_valid),
    .io_reservationStation_bits_destinationTag_threadId(executors_1_io_reservationStation_bits_destinationTag_threadId),
    .io_reservationStation_bits_destinationTag_id(executors_1_io_reservationStation_bits_destinationTag_id),
    .io_reservationStation_bits_value1(executors_1_io_reservationStation_bits_value1),
    .io_reservationStation_bits_value2(executors_1_io_reservationStation_bits_value2),
    .io_reservationStation_bits_function3(executors_1_io_reservationStation_bits_function3),
    .io_reservationStation_bits_immediateOrFunction7(executors_1_io_reservationStation_bits_immediateOrFunction7),
    .io_reservationStation_bits_opcode(executors_1_io_reservationStation_bits_opcode),
    .io_reservationStation_bits_wasCompressed(executors_1_io_reservationStation_bits_wasCompressed),
    .io_out_ready(executors_1_io_out_ready),
    .io_out_valid(executors_1_io_out_valid),
    .io_out_bits_resultType(executors_1_io_out_bits_resultType),
    .io_out_bits_value(executors_1_io_out_bits_value),
    .io_out_bits_tag_threadId(executors_1_io_out_bits_tag_threadId),
    .io_out_bits_tag_id(executors_1_io_out_bits_tag_id),
    .io_fetch_ready(executors_1_io_fetch_ready),
    .io_fetch_valid(executors_1_io_fetch_valid),
    .io_fetch_bits_threadId(executors_1_io_fetch_bits_threadId),
    .io_fetch_bits_programCounterOffset(executors_1_io_fetch_bits_programCounterOffset)
  );
  ExternalMemoryInterface externalMemoryInterface ( // @[B4Processor.scala 59:47]
    .clock(externalMemoryInterface_clock),
    .reset(externalMemoryInterface_reset),
    .io_dataWriteRequests_ready(externalMemoryInterface_io_dataWriteRequests_ready),
    .io_dataWriteRequests_valid(externalMemoryInterface_io_dataWriteRequests_valid),
    .io_dataWriteRequests_bits_address(externalMemoryInterface_io_dataWriteRequests_bits_address),
    .io_dataWriteRequests_bits_data(externalMemoryInterface_io_dataWriteRequests_bits_data),
    .io_dataWriteRequests_bits_mask(externalMemoryInterface_io_dataWriteRequests_bits_mask),
    .io_dataReadRequests_ready(externalMemoryInterface_io_dataReadRequests_ready),
    .io_dataReadRequests_valid(externalMemoryInterface_io_dataReadRequests_valid),
    .io_dataReadRequests_bits_address(externalMemoryInterface_io_dataReadRequests_bits_address),
    .io_dataReadRequests_bits_size(externalMemoryInterface_io_dataReadRequests_bits_size),
    .io_dataReadRequests_bits_signed(externalMemoryInterface_io_dataReadRequests_bits_signed),
    .io_dataReadRequests_bits_outputTag_threadId(externalMemoryInterface_io_dataReadRequests_bits_outputTag_threadId),
    .io_dataReadRequests_bits_outputTag_id(externalMemoryInterface_io_dataReadRequests_bits_outputTag_id),
    .io_instructionFetchRequest_0_ready(externalMemoryInterface_io_instructionFetchRequest_0_ready),
    .io_instructionFetchRequest_0_valid(externalMemoryInterface_io_instructionFetchRequest_0_valid),
    .io_instructionFetchRequest_0_bits_address(externalMemoryInterface_io_instructionFetchRequest_0_bits_address),
    .io_instructionFetchRequest_1_ready(externalMemoryInterface_io_instructionFetchRequest_1_ready),
    .io_instructionFetchRequest_1_valid(externalMemoryInterface_io_instructionFetchRequest_1_valid),
    .io_instructionFetchRequest_1_bits_address(externalMemoryInterface_io_instructionFetchRequest_1_bits_address),
    .io_dataReadOut_ready(externalMemoryInterface_io_dataReadOut_ready),
    .io_dataReadOut_valid(externalMemoryInterface_io_dataReadOut_valid),
    .io_dataReadOut_bits_value(externalMemoryInterface_io_dataReadOut_bits_value),
    .io_dataReadOut_bits_isError(externalMemoryInterface_io_dataReadOut_bits_isError),
    .io_dataReadOut_bits_tag_threadId(externalMemoryInterface_io_dataReadOut_bits_tag_threadId),
    .io_dataReadOut_bits_tag_id(externalMemoryInterface_io_dataReadOut_bits_tag_id),
    .io_instructionOut_0_valid(externalMemoryInterface_io_instructionOut_0_valid),
    .io_instructionOut_0_bits_inner(externalMemoryInterface_io_instructionOut_0_bits_inner),
    .io_instructionOut_1_valid(externalMemoryInterface_io_instructionOut_1_valid),
    .io_instructionOut_1_bits_inner(externalMemoryInterface_io_instructionOut_1_bits_inner),
    .io_coordinator_writeAddress_ready(externalMemoryInterface_io_coordinator_writeAddress_ready),
    .io_coordinator_writeAddress_valid(externalMemoryInterface_io_coordinator_writeAddress_valid),
    .io_coordinator_writeAddress_bits_ADDR(externalMemoryInterface_io_coordinator_writeAddress_bits_ADDR),
    .io_coordinator_writeAddress_bits_CACHE(externalMemoryInterface_io_coordinator_writeAddress_bits_CACHE),
    .io_coordinator_write_ready(externalMemoryInterface_io_coordinator_write_ready),
    .io_coordinator_write_valid(externalMemoryInterface_io_coordinator_write_valid),
    .io_coordinator_write_bits_DATA(externalMemoryInterface_io_coordinator_write_bits_DATA),
    .io_coordinator_write_bits_STRB(externalMemoryInterface_io_coordinator_write_bits_STRB),
    .io_coordinator_write_bits_LAST(externalMemoryInterface_io_coordinator_write_bits_LAST),
    .io_coordinator_writeResponse_ready(externalMemoryInterface_io_coordinator_writeResponse_ready),
    .io_coordinator_writeResponse_valid(externalMemoryInterface_io_coordinator_writeResponse_valid),
    .io_coordinator_readAddress_ready(externalMemoryInterface_io_coordinator_readAddress_ready),
    .io_coordinator_readAddress_valid(externalMemoryInterface_io_coordinator_readAddress_valid),
    .io_coordinator_readAddress_bits_ADDR(externalMemoryInterface_io_coordinator_readAddress_bits_ADDR),
    .io_coordinator_readAddress_bits_LEN(externalMemoryInterface_io_coordinator_readAddress_bits_LEN),
    .io_coordinator_readAddress_bits_CACHE(externalMemoryInterface_io_coordinator_readAddress_bits_CACHE),
    .io_coordinator_read_ready(externalMemoryInterface_io_coordinator_read_ready),
    .io_coordinator_read_valid(externalMemoryInterface_io_coordinator_read_valid),
    .io_coordinator_read_bits_DATA(externalMemoryInterface_io_coordinator_read_bits_DATA),
    .io_coordinator_read_bits_RESP(externalMemoryInterface_io_coordinator_read_bits_RESP)
  );
  CSRReservationStation csrReservationStation_0 ( // @[B4Processor.scala 62:36]
    .clock(csrReservationStation_0_clock),
    .reset(csrReservationStation_0_reset),
    .io_decoderInput_0_ready(csrReservationStation_0_io_decoderInput_0_ready),
    .io_decoderInput_0_valid(csrReservationStation_0_io_decoderInput_0_valid),
    .io_decoderInput_0_bits_sourceTag_threadId(csrReservationStation_0_io_decoderInput_0_bits_sourceTag_threadId),
    .io_decoderInput_0_bits_sourceTag_id(csrReservationStation_0_io_decoderInput_0_bits_sourceTag_id),
    .io_decoderInput_0_bits_destinationTag_threadId(
      csrReservationStation_0_io_decoderInput_0_bits_destinationTag_threadId),
    .io_decoderInput_0_bits_destinationTag_id(csrReservationStation_0_io_decoderInput_0_bits_destinationTag_id),
    .io_decoderInput_0_bits_value(csrReservationStation_0_io_decoderInput_0_bits_value),
    .io_decoderInput_0_bits_ready(csrReservationStation_0_io_decoderInput_0_bits_ready),
    .io_decoderInput_0_bits_address(csrReservationStation_0_io_decoderInput_0_bits_address),
    .io_decoderInput_0_bits_csrAccessType(csrReservationStation_0_io_decoderInput_0_bits_csrAccessType),
    .io_toCSR_ready(csrReservationStation_0_io_toCSR_ready),
    .io_toCSR_valid(csrReservationStation_0_io_toCSR_valid),
    .io_toCSR_bits_address(csrReservationStation_0_io_toCSR_bits_address),
    .io_toCSR_bits_value(csrReservationStation_0_io_toCSR_bits_value),
    .io_toCSR_bits_destinationTag_threadId(csrReservationStation_0_io_toCSR_bits_destinationTag_threadId),
    .io_toCSR_bits_destinationTag_id(csrReservationStation_0_io_toCSR_bits_destinationTag_id),
    .io_toCSR_bits_csrAccessType(csrReservationStation_0_io_toCSR_bits_csrAccessType),
    .io_output_outputs_valid(csrReservationStation_0_io_output_outputs_valid),
    .io_output_outputs_bits_value(csrReservationStation_0_io_output_outputs_bits_value),
    .io_output_outputs_bits_tag_threadId(csrReservationStation_0_io_output_outputs_bits_tag_threadId),
    .io_output_outputs_bits_tag_id(csrReservationStation_0_io_output_outputs_bits_tag_id),
    .io_empty(csrReservationStation_0_io_empty)
  );
  CSRReservationStation csrReservationStation_1 ( // @[B4Processor.scala 62:36]
    .clock(csrReservationStation_1_clock),
    .reset(csrReservationStation_1_reset),
    .io_decoderInput_0_ready(csrReservationStation_1_io_decoderInput_0_ready),
    .io_decoderInput_0_valid(csrReservationStation_1_io_decoderInput_0_valid),
    .io_decoderInput_0_bits_sourceTag_threadId(csrReservationStation_1_io_decoderInput_0_bits_sourceTag_threadId),
    .io_decoderInput_0_bits_sourceTag_id(csrReservationStation_1_io_decoderInput_0_bits_sourceTag_id),
    .io_decoderInput_0_bits_destinationTag_threadId(
      csrReservationStation_1_io_decoderInput_0_bits_destinationTag_threadId),
    .io_decoderInput_0_bits_destinationTag_id(csrReservationStation_1_io_decoderInput_0_bits_destinationTag_id),
    .io_decoderInput_0_bits_value(csrReservationStation_1_io_decoderInput_0_bits_value),
    .io_decoderInput_0_bits_ready(csrReservationStation_1_io_decoderInput_0_bits_ready),
    .io_decoderInput_0_bits_address(csrReservationStation_1_io_decoderInput_0_bits_address),
    .io_decoderInput_0_bits_csrAccessType(csrReservationStation_1_io_decoderInput_0_bits_csrAccessType),
    .io_toCSR_ready(csrReservationStation_1_io_toCSR_ready),
    .io_toCSR_valid(csrReservationStation_1_io_toCSR_valid),
    .io_toCSR_bits_address(csrReservationStation_1_io_toCSR_bits_address),
    .io_toCSR_bits_value(csrReservationStation_1_io_toCSR_bits_value),
    .io_toCSR_bits_destinationTag_threadId(csrReservationStation_1_io_toCSR_bits_destinationTag_threadId),
    .io_toCSR_bits_destinationTag_id(csrReservationStation_1_io_toCSR_bits_destinationTag_id),
    .io_toCSR_bits_csrAccessType(csrReservationStation_1_io_toCSR_bits_csrAccessType),
    .io_output_outputs_valid(csrReservationStation_1_io_output_outputs_valid),
    .io_output_outputs_bits_value(csrReservationStation_1_io_output_outputs_bits_value),
    .io_output_outputs_bits_tag_threadId(csrReservationStation_1_io_output_outputs_bits_tag_threadId),
    .io_output_outputs_bits_tag_id(csrReservationStation_1_io_output_outputs_bits_tag_id),
    .io_empty(csrReservationStation_1_io_empty)
  );
  CSR csr_0 ( // @[B4Processor.scala 63:61]
    .clock(csr_0_clock),
    .reset(csr_0_reset),
    .io_decoderInput_ready(csr_0_io_decoderInput_ready),
    .io_decoderInput_valid(csr_0_io_decoderInput_valid),
    .io_decoderInput_bits_address(csr_0_io_decoderInput_bits_address),
    .io_decoderInput_bits_value(csr_0_io_decoderInput_bits_value),
    .io_decoderInput_bits_destinationTag_threadId(csr_0_io_decoderInput_bits_destinationTag_threadId),
    .io_decoderInput_bits_destinationTag_id(csr_0_io_decoderInput_bits_destinationTag_id),
    .io_decoderInput_bits_csrAccessType(csr_0_io_decoderInput_bits_csrAccessType),
    .io_CSROutput_ready(csr_0_io_CSROutput_ready),
    .io_CSROutput_valid(csr_0_io_CSROutput_valid),
    .io_CSROutput_bits_value(csr_0_io_CSROutput_bits_value),
    .io_CSROutput_bits_isError(csr_0_io_CSROutput_bits_isError),
    .io_CSROutput_bits_tag_threadId(csr_0_io_CSROutput_bits_tag_threadId),
    .io_CSROutput_bits_tag_id(csr_0_io_CSROutput_bits_tag_id),
    .io_fetch_mtvec(csr_0_io_fetch_mtvec),
    .io_fetch_mepc(csr_0_io_fetch_mepc),
    .io_fetch_mcause(csr_0_io_fetch_mcause),
    .io_reorderBuffer_retireCount(csr_0_io_reorderBuffer_retireCount)
  );
  CSR_1 csr_1 ( // @[B4Processor.scala 63:61]
    .clock(csr_1_clock),
    .reset(csr_1_reset),
    .io_decoderInput_ready(csr_1_io_decoderInput_ready),
    .io_decoderInput_valid(csr_1_io_decoderInput_valid),
    .io_decoderInput_bits_address(csr_1_io_decoderInput_bits_address),
    .io_decoderInput_bits_value(csr_1_io_decoderInput_bits_value),
    .io_decoderInput_bits_destinationTag_threadId(csr_1_io_decoderInput_bits_destinationTag_threadId),
    .io_decoderInput_bits_destinationTag_id(csr_1_io_decoderInput_bits_destinationTag_id),
    .io_decoderInput_bits_csrAccessType(csr_1_io_decoderInput_bits_csrAccessType),
    .io_CSROutput_ready(csr_1_io_CSROutput_ready),
    .io_CSROutput_valid(csr_1_io_CSROutput_valid),
    .io_CSROutput_bits_value(csr_1_io_CSROutput_bits_value),
    .io_CSROutput_bits_isError(csr_1_io_CSROutput_bits_isError),
    .io_CSROutput_bits_tag_threadId(csr_1_io_CSROutput_bits_tag_threadId),
    .io_CSROutput_bits_tag_id(csr_1_io_CSROutput_bits_tag_id),
    .io_fetch_mtvec(csr_1_io_fetch_mtvec),
    .io_fetch_mepc(csr_1_io_fetch_mepc),
    .io_fetch_mcause(csr_1_io_fetch_mcause),
    .io_reorderBuffer_retireCount(csr_1_io_reorderBuffer_retireCount)
  );
  assign axi_writeAddress_valid = externalMemoryInterface_io_coordinator_writeAddress_valid; // @[B4Processor.scala 65:7]
  assign axi_writeAddress_bits_ADDR = externalMemoryInterface_io_coordinator_writeAddress_bits_ADDR; // @[B4Processor.scala 65:7]
  assign axi_writeAddress_bits_LEN = 8'h0; // @[B4Processor.scala 65:7]
  assign axi_writeAddress_bits_SIZE = 3'h6; // @[B4Processor.scala 65:7]
  assign axi_writeAddress_bits_BURST = 2'h1; // @[B4Processor.scala 65:7]
  assign axi_writeAddress_bits_LOCK = 1'h0; // @[B4Processor.scala 65:7]
  assign axi_writeAddress_bits_CACHE = externalMemoryInterface_io_coordinator_writeAddress_bits_CACHE; // @[B4Processor.scala 65:7]
  assign axi_writeAddress_bits_PROT = 3'h0; // @[B4Processor.scala 65:7]
  assign axi_writeAddress_bits_QOS = 4'h0; // @[B4Processor.scala 65:7]
  assign axi_writeAddress_bits_REGION = 4'h0; // @[B4Processor.scala 65:7]
  assign axi_write_valid = externalMemoryInterface_io_coordinator_write_valid; // @[B4Processor.scala 65:7]
  assign axi_write_bits_DATA = externalMemoryInterface_io_coordinator_write_bits_DATA; // @[B4Processor.scala 65:7]
  assign axi_write_bits_STRB = externalMemoryInterface_io_coordinator_write_bits_STRB; // @[B4Processor.scala 65:7]
  assign axi_write_bits_LAST = externalMemoryInterface_io_coordinator_write_bits_LAST; // @[B4Processor.scala 65:7]
  assign axi_writeResponse_ready = externalMemoryInterface_io_coordinator_writeResponse_ready; // @[B4Processor.scala 65:7]
  assign axi_readAddress_valid = externalMemoryInterface_io_coordinator_readAddress_valid; // @[B4Processor.scala 65:7]
  assign axi_readAddress_bits_ADDR = externalMemoryInterface_io_coordinator_readAddress_bits_ADDR; // @[B4Processor.scala 65:7]
  assign axi_readAddress_bits_LEN = externalMemoryInterface_io_coordinator_readAddress_bits_LEN; // @[B4Processor.scala 65:7]
  assign axi_readAddress_bits_SIZE = 3'h6; // @[B4Processor.scala 65:7]
  assign axi_readAddress_bits_BURST = 2'h1; // @[B4Processor.scala 65:7]
  assign axi_readAddress_bits_LOCK = 1'h0; // @[B4Processor.scala 65:7]
  assign axi_readAddress_bits_CACHE = externalMemoryInterface_io_coordinator_readAddress_bits_CACHE; // @[B4Processor.scala 65:7]
  assign axi_readAddress_bits_PROT = 3'h0; // @[B4Processor.scala 65:7]
  assign axi_readAddress_bits_QOS = 4'h0; // @[B4Processor.scala 65:7]
  assign axi_readAddress_bits_REGION = 4'h0; // @[B4Processor.scala 65:7]
  assign axi_read_ready = externalMemoryInterface_io_coordinator_read_ready; // @[B4Processor.scala 65:7]
  assign instructionCache_0_clock = clock;
  assign instructionCache_0_reset = reset;
  assign instructionCache_0_io_fetch_0_address_valid = fetch_0_io_cache_0_address_valid; // @[B4Processor.scala 101:36]
  assign instructionCache_0_io_fetch_0_address_bits = fetch_0_io_cache_0_address_bits; // @[B4Processor.scala 101:36]
  assign instructionCache_0_io_memory_request_ready = externalMemoryInterface_io_instructionFetchRequest_0_ready; // @[B4Processor.scala 178:61]
  assign instructionCache_0_io_memory_response_valid = externalMemoryInterface_io_instructionOut_0_valid; // @[B4Processor.scala 181:52]
  assign instructionCache_0_io_memory_response_bits_inner = externalMemoryInterface_io_instructionOut_0_bits_inner; // @[B4Processor.scala 181:52]
  assign instructionCache_1_clock = clock;
  assign instructionCache_1_reset = reset;
  assign instructionCache_1_io_fetch_0_address_valid = fetch_1_io_cache_0_address_valid; // @[B4Processor.scala 101:36]
  assign instructionCache_1_io_fetch_0_address_bits = fetch_1_io_cache_0_address_bits; // @[B4Processor.scala 101:36]
  assign instructionCache_1_io_memory_request_ready = externalMemoryInterface_io_instructionFetchRequest_1_ready; // @[B4Processor.scala 178:61]
  assign instructionCache_1_io_memory_response_valid = externalMemoryInterface_io_instructionOut_1_valid; // @[B4Processor.scala 181:52]
  assign instructionCache_1_io_memory_response_bits_inner = externalMemoryInterface_io_instructionOut_1_bits_inner; // @[B4Processor.scala 181:52]
  assign fetch_0_clock = clock;
  assign fetch_0_reset = reset;
  assign fetch_0_io_cache_0_output_valid = instructionCache_0_io_fetch_0_output_valid; // @[B4Processor.scala 101:36]
  assign fetch_0_io_cache_0_output_bits = instructionCache_0_io_fetch_0_output_bits; // @[B4Processor.scala 101:36]
  assign fetch_0_io_reorderBufferEmpty = reorderBuffer_0_io_isEmpty; // @[B4Processor.scala 166:38]
  assign fetch_0_io_loadStoreQueueEmpty = loadStoreQueue_0_io_isEmpty; // @[B4Processor.scala 163:39]
  assign fetch_0_io_collectedBranchAddresses_addresses_valid = branchAddressCollector_io_fetch_0_addresses_valid; // @[B4Processor.scala 153:44]
  assign fetch_0_io_collectedBranchAddresses_addresses_bits_threadId =
    branchAddressCollector_io_fetch_0_addresses_bits_threadId; // @[B4Processor.scala 153:44]
  assign fetch_0_io_collectedBranchAddresses_addresses_bits_programCounterOffset =
    branchAddressCollector_io_fetch_0_addresses_bits_programCounterOffset; // @[B4Processor.scala 153:44]
  assign fetch_0_io_fetchBuffer_toBuffer_0_ready = fetchBuffer_0_io_input_toBuffer_0_ready; // @[B4Processor.scala 104:31]
  assign fetch_0_io_fetchBuffer_empty = fetchBuffer_0_io_input_empty; // @[B4Processor.scala 104:31]
  assign fetch_0_io_csr_mtvec = csr_0_io_fetch_mtvec; // @[B4Processor.scala 114:23]
  assign fetch_0_io_csr_mepc = csr_0_io_fetch_mepc; // @[B4Processor.scala 114:23]
  assign fetch_0_io_csr_mcause = csr_0_io_fetch_mcause; // @[B4Processor.scala 114:23]
  assign fetch_0_io_csrReservationStationEmpty = csrReservationStation_0_io_empty; // @[B4Processor.scala 116:46]
  assign fetch_0_io_isError = reorderBuffer_0_io_isError; // @[B4Processor.scala 121:27]
  assign fetch_1_clock = clock;
  assign fetch_1_reset = reset;
  assign fetch_1_io_cache_0_output_valid = instructionCache_1_io_fetch_0_output_valid; // @[B4Processor.scala 101:36]
  assign fetch_1_io_cache_0_output_bits = instructionCache_1_io_fetch_0_output_bits; // @[B4Processor.scala 101:36]
  assign fetch_1_io_reorderBufferEmpty = reorderBuffer_1_io_isEmpty; // @[B4Processor.scala 166:38]
  assign fetch_1_io_loadStoreQueueEmpty = loadStoreQueue_1_io_isEmpty; // @[B4Processor.scala 163:39]
  assign fetch_1_io_collectedBranchAddresses_addresses_valid = branchAddressCollector_io_fetch_1_addresses_valid; // @[B4Processor.scala 153:44]
  assign fetch_1_io_collectedBranchAddresses_addresses_bits_threadId =
    branchAddressCollector_io_fetch_1_addresses_bits_threadId; // @[B4Processor.scala 153:44]
  assign fetch_1_io_collectedBranchAddresses_addresses_bits_programCounterOffset =
    branchAddressCollector_io_fetch_1_addresses_bits_programCounterOffset; // @[B4Processor.scala 153:44]
  assign fetch_1_io_fetchBuffer_toBuffer_0_ready = fetchBuffer_1_io_input_toBuffer_0_ready; // @[B4Processor.scala 104:31]
  assign fetch_1_io_fetchBuffer_empty = fetchBuffer_1_io_input_empty; // @[B4Processor.scala 104:31]
  assign fetch_1_io_csr_mtvec = csr_1_io_fetch_mtvec; // @[B4Processor.scala 114:23]
  assign fetch_1_io_csr_mepc = csr_1_io_fetch_mepc; // @[B4Processor.scala 114:23]
  assign fetch_1_io_csr_mcause = csr_1_io_fetch_mcause; // @[B4Processor.scala 114:23]
  assign fetch_1_io_csrReservationStationEmpty = csrReservationStation_1_io_empty; // @[B4Processor.scala 116:46]
  assign fetch_1_io_isError = reorderBuffer_1_io_isError; // @[B4Processor.scala 121:27]
  assign fetchBuffer_0_clock = clock;
  assign fetchBuffer_0_reset = reset;
  assign fetchBuffer_0_io_output_0_ready = uncompresser_0_0_io_fetch_ready; // @[B4Processor.scala 127:37]
  assign fetchBuffer_0_io_input_toBuffer_0_valid = fetch_0_io_fetchBuffer_toBuffer_0_valid; // @[B4Processor.scala 104:31]
  assign fetchBuffer_0_io_input_toBuffer_0_bits_instruction = fetch_0_io_fetchBuffer_toBuffer_0_bits_instruction; // @[B4Processor.scala 104:31]
  assign fetchBuffer_0_io_input_toBuffer_0_bits_programCounter = fetch_0_io_fetchBuffer_toBuffer_0_bits_programCounter; // @[B4Processor.scala 104:31]
  assign fetchBuffer_1_clock = clock;
  assign fetchBuffer_1_reset = reset;
  assign fetchBuffer_1_io_output_0_ready = uncompresser_1_0_io_fetch_ready; // @[B4Processor.scala 127:37]
  assign fetchBuffer_1_io_input_toBuffer_0_valid = fetch_1_io_fetchBuffer_toBuffer_0_valid; // @[B4Processor.scala 104:31]
  assign fetchBuffer_1_io_input_toBuffer_0_bits_instruction = fetch_1_io_fetchBuffer_toBuffer_0_bits_instruction; // @[B4Processor.scala 104:31]
  assign fetchBuffer_1_io_input_toBuffer_0_bits_programCounter = fetch_1_io_fetchBuffer_toBuffer_0_bits_programCounter; // @[B4Processor.scala 104:31]
  assign reorderBuffer_0_clock = clock;
  assign reorderBuffer_0_reset = reset;
  assign reorderBuffer_0_io_decoders_0_source1_sourceRegister = decoders_0_0_io_reorderBuffer_source1_sourceRegister; // @[B4Processor.scala 133:41]
  assign reorderBuffer_0_io_decoders_0_source2_sourceRegister = decoders_0_0_io_reorderBuffer_source2_sourceRegister; // @[B4Processor.scala 133:41]
  assign reorderBuffer_0_io_decoders_0_destination_destinationRegister =
    decoders_0_0_io_reorderBuffer_destination_destinationRegister; // @[B4Processor.scala 133:41]
  assign reorderBuffer_0_io_decoders_0_destination_storeSign = decoders_0_0_io_reorderBuffer_destination_storeSign; // @[B4Processor.scala 133:41]
  assign reorderBuffer_0_io_decoders_0_valid = decoders_0_0_io_reorderBuffer_valid; // @[B4Processor.scala 133:41]
  assign reorderBuffer_0_io_collectedOutputs_outputs_valid = outputCollector_io_outputs_0_outputs_valid; // @[B4Processor.scala 172:44]
  assign reorderBuffer_0_io_collectedOutputs_outputs_bits_resultType =
    outputCollector_io_outputs_0_outputs_bits_resultType; // @[B4Processor.scala 172:44]
  assign reorderBuffer_0_io_collectedOutputs_outputs_bits_value = outputCollector_io_outputs_0_outputs_bits_value; // @[B4Processor.scala 172:44]
  assign reorderBuffer_0_io_collectedOutputs_outputs_bits_isError = outputCollector_io_outputs_0_outputs_bits_isError; // @[B4Processor.scala 172:44]
  assign reorderBuffer_0_io_collectedOutputs_outputs_bits_tag_threadId =
    outputCollector_io_outputs_0_outputs_bits_tag_threadId; // @[B4Processor.scala 172:44]
  assign reorderBuffer_0_io_collectedOutputs_outputs_bits_tag_id = outputCollector_io_outputs_0_outputs_bits_tag_id; // @[B4Processor.scala 172:44]
  assign reorderBuffer_1_clock = clock;
  assign reorderBuffer_1_reset = reset;
  assign reorderBuffer_1_io_decoders_0_source1_sourceRegister = decoders_1_0_io_reorderBuffer_source1_sourceRegister; // @[B4Processor.scala 133:41]
  assign reorderBuffer_1_io_decoders_0_source2_sourceRegister = decoders_1_0_io_reorderBuffer_source2_sourceRegister; // @[B4Processor.scala 133:41]
  assign reorderBuffer_1_io_decoders_0_destination_destinationRegister =
    decoders_1_0_io_reorderBuffer_destination_destinationRegister; // @[B4Processor.scala 133:41]
  assign reorderBuffer_1_io_decoders_0_destination_storeSign = decoders_1_0_io_reorderBuffer_destination_storeSign; // @[B4Processor.scala 133:41]
  assign reorderBuffer_1_io_decoders_0_valid = decoders_1_0_io_reorderBuffer_valid; // @[B4Processor.scala 133:41]
  assign reorderBuffer_1_io_collectedOutputs_outputs_valid = outputCollector_io_outputs_1_outputs_valid; // @[B4Processor.scala 172:44]
  assign reorderBuffer_1_io_collectedOutputs_outputs_bits_resultType =
    outputCollector_io_outputs_1_outputs_bits_resultType; // @[B4Processor.scala 172:44]
  assign reorderBuffer_1_io_collectedOutputs_outputs_bits_value = outputCollector_io_outputs_1_outputs_bits_value; // @[B4Processor.scala 172:44]
  assign reorderBuffer_1_io_collectedOutputs_outputs_bits_isError = outputCollector_io_outputs_1_outputs_bits_isError; // @[B4Processor.scala 172:44]
  assign reorderBuffer_1_io_collectedOutputs_outputs_bits_tag_threadId =
    outputCollector_io_outputs_1_outputs_bits_tag_threadId; // @[B4Processor.scala 172:44]
  assign reorderBuffer_1_io_collectedOutputs_outputs_bits_tag_id = outputCollector_io_outputs_1_outputs_bits_tag_id; // @[B4Processor.scala 172:44]
  assign registerFile_0_clock = clock;
  assign registerFile_0_reset = reset;
  assign registerFile_0_io_decoders_0_sourceRegister1 = decoders_0_0_io_registerFile_sourceRegister1; // @[B4Processor.scala 140:40]
  assign registerFile_0_io_decoders_0_sourceRegister2 = decoders_0_0_io_registerFile_sourceRegister2; // @[B4Processor.scala 140:40]
  assign registerFile_0_io_reorderBuffer_0_valid = reorderBuffer_0_io_registerFile_0_valid; // @[B4Processor.scala 160:40]
  assign registerFile_0_io_reorderBuffer_0_bits_destinationRegister =
    reorderBuffer_0_io_registerFile_0_bits_destinationRegister; // @[B4Processor.scala 160:40]
  assign registerFile_0_io_reorderBuffer_0_bits_value = reorderBuffer_0_io_registerFile_0_bits_value; // @[B4Processor.scala 160:40]
  assign registerFile_0_io_reorderBuffer_1_valid = reorderBuffer_0_io_registerFile_1_valid; // @[B4Processor.scala 160:40]
  assign registerFile_0_io_reorderBuffer_1_bits_destinationRegister =
    reorderBuffer_0_io_registerFile_1_bits_destinationRegister; // @[B4Processor.scala 160:40]
  assign registerFile_0_io_reorderBuffer_1_bits_value = reorderBuffer_0_io_registerFile_1_bits_value; // @[B4Processor.scala 160:40]
  assign registerFile_0_io_reorderBuffer_2_valid = reorderBuffer_0_io_registerFile_2_valid; // @[B4Processor.scala 160:40]
  assign registerFile_0_io_reorderBuffer_2_bits_destinationRegister =
    reorderBuffer_0_io_registerFile_2_bits_destinationRegister; // @[B4Processor.scala 160:40]
  assign registerFile_0_io_reorderBuffer_2_bits_value = reorderBuffer_0_io_registerFile_2_bits_value; // @[B4Processor.scala 160:40]
  assign registerFile_0_io_reorderBuffer_3_valid = reorderBuffer_0_io_registerFile_3_valid; // @[B4Processor.scala 160:40]
  assign registerFile_0_io_reorderBuffer_3_bits_destinationRegister =
    reorderBuffer_0_io_registerFile_3_bits_destinationRegister; // @[B4Processor.scala 160:40]
  assign registerFile_0_io_reorderBuffer_3_bits_value = reorderBuffer_0_io_registerFile_3_bits_value; // @[B4Processor.scala 160:40]
  assign registerFile_1_clock = clock;
  assign registerFile_1_reset = reset;
  assign registerFile_1_io_decoders_0_sourceRegister1 = decoders_1_0_io_registerFile_sourceRegister1; // @[B4Processor.scala 140:40]
  assign registerFile_1_io_decoders_0_sourceRegister2 = decoders_1_0_io_registerFile_sourceRegister2; // @[B4Processor.scala 140:40]
  assign registerFile_1_io_reorderBuffer_0_valid = reorderBuffer_1_io_registerFile_0_valid; // @[B4Processor.scala 160:40]
  assign registerFile_1_io_reorderBuffer_0_bits_destinationRegister =
    reorderBuffer_1_io_registerFile_0_bits_destinationRegister; // @[B4Processor.scala 160:40]
  assign registerFile_1_io_reorderBuffer_0_bits_value = reorderBuffer_1_io_registerFile_0_bits_value; // @[B4Processor.scala 160:40]
  assign registerFile_1_io_reorderBuffer_1_valid = reorderBuffer_1_io_registerFile_1_valid; // @[B4Processor.scala 160:40]
  assign registerFile_1_io_reorderBuffer_1_bits_destinationRegister =
    reorderBuffer_1_io_registerFile_1_bits_destinationRegister; // @[B4Processor.scala 160:40]
  assign registerFile_1_io_reorderBuffer_1_bits_value = reorderBuffer_1_io_registerFile_1_bits_value; // @[B4Processor.scala 160:40]
  assign registerFile_1_io_reorderBuffer_2_valid = reorderBuffer_1_io_registerFile_2_valid; // @[B4Processor.scala 160:40]
  assign registerFile_1_io_reorderBuffer_2_bits_destinationRegister =
    reorderBuffer_1_io_registerFile_2_bits_destinationRegister; // @[B4Processor.scala 160:40]
  assign registerFile_1_io_reorderBuffer_2_bits_value = reorderBuffer_1_io_registerFile_2_bits_value; // @[B4Processor.scala 160:40]
  assign registerFile_1_io_reorderBuffer_3_valid = reorderBuffer_1_io_registerFile_3_valid; // @[B4Processor.scala 160:40]
  assign registerFile_1_io_reorderBuffer_3_bits_destinationRegister =
    reorderBuffer_1_io_registerFile_3_bits_destinationRegister; // @[B4Processor.scala 160:40]
  assign registerFile_1_io_reorderBuffer_3_bits_value = reorderBuffer_1_io_registerFile_3_bits_value; // @[B4Processor.scala 160:40]
  assign loadStoreQueue_0_clock = clock;
  assign loadStoreQueue_0_reset = reset;
  assign loadStoreQueue_0_io_decoders_0_valid = decoders_0_0_io_loadStoreQueue_valid; // @[B4Processor.scala 149:42]
  assign loadStoreQueue_0_io_decoders_0_bits_accessInfo_accessType =
    decoders_0_0_io_loadStoreQueue_bits_accessInfo_accessType; // @[B4Processor.scala 149:42]
  assign loadStoreQueue_0_io_decoders_0_bits_accessInfo_signed = decoders_0_0_io_loadStoreQueue_bits_accessInfo_signed; // @[B4Processor.scala 149:42]
  assign loadStoreQueue_0_io_decoders_0_bits_accessInfo_accessWidth =
    decoders_0_0_io_loadStoreQueue_bits_accessInfo_accessWidth; // @[B4Processor.scala 149:42]
  assign loadStoreQueue_0_io_decoders_0_bits_addressAndLoadResultTag_threadId =
    decoders_0_0_io_loadStoreQueue_bits_addressAndLoadResultTag_threadId; // @[B4Processor.scala 149:42]
  assign loadStoreQueue_0_io_decoders_0_bits_addressAndLoadResultTag_id =
    decoders_0_0_io_loadStoreQueue_bits_addressAndLoadResultTag_id; // @[B4Processor.scala 149:42]
  assign loadStoreQueue_0_io_decoders_0_bits_address = decoders_0_0_io_loadStoreQueue_bits_address; // @[B4Processor.scala 149:42]
  assign loadStoreQueue_0_io_decoders_0_bits_addressValid = decoders_0_0_io_loadStoreQueue_bits_addressValid; // @[B4Processor.scala 149:42]
  assign loadStoreQueue_0_io_decoders_0_bits_storeDataTag_threadId =
    decoders_0_0_io_loadStoreQueue_bits_storeDataTag_threadId; // @[B4Processor.scala 149:42]
  assign loadStoreQueue_0_io_decoders_0_bits_storeDataTag_id = decoders_0_0_io_loadStoreQueue_bits_storeDataTag_id; // @[B4Processor.scala 149:42]
  assign loadStoreQueue_0_io_decoders_0_bits_storeData = decoders_0_0_io_loadStoreQueue_bits_storeData; // @[B4Processor.scala 149:42]
  assign loadStoreQueue_0_io_decoders_0_bits_storeDataValid = decoders_0_0_io_loadStoreQueue_bits_storeDataValid; // @[B4Processor.scala 149:42]
  assign loadStoreQueue_0_io_outputCollector_outputs_valid = outputCollector_io_outputs_0_outputs_valid; // @[B4Processor.scala 157:44]
  assign loadStoreQueue_0_io_outputCollector_outputs_bits_resultType =
    outputCollector_io_outputs_0_outputs_bits_resultType; // @[B4Processor.scala 157:44]
  assign loadStoreQueue_0_io_outputCollector_outputs_bits_value = outputCollector_io_outputs_0_outputs_bits_value; // @[B4Processor.scala 157:44]
  assign loadStoreQueue_0_io_outputCollector_outputs_bits_tag_threadId =
    outputCollector_io_outputs_0_outputs_bits_tag_threadId; // @[B4Processor.scala 157:44]
  assign loadStoreQueue_0_io_outputCollector_outputs_bits_tag_id = outputCollector_io_outputs_0_outputs_bits_tag_id; // @[B4Processor.scala 157:44]
  assign loadStoreQueue_0_io_reorderBuffer_0_valid = reorderBuffer_0_io_loadStoreQueue_0_valid; // @[B4Processor.scala 175:42]
  assign loadStoreQueue_0_io_reorderBuffer_0_bits_destinationTag_threadId = 1'h0; // @[B4Processor.scala 175:42]
  assign loadStoreQueue_0_io_reorderBuffer_0_bits_destinationTag_id =
    reorderBuffer_0_io_loadStoreQueue_0_bits_destinationTag_id; // @[B4Processor.scala 175:42]
  assign loadStoreQueue_0_io_reorderBuffer_1_valid = reorderBuffer_0_io_loadStoreQueue_1_valid; // @[B4Processor.scala 175:42]
  assign loadStoreQueue_0_io_reorderBuffer_1_bits_destinationTag_threadId = 1'h0; // @[B4Processor.scala 175:42]
  assign loadStoreQueue_0_io_reorderBuffer_1_bits_destinationTag_id =
    reorderBuffer_0_io_loadStoreQueue_1_bits_destinationTag_id; // @[B4Processor.scala 175:42]
  assign loadStoreQueue_0_io_reorderBuffer_2_valid = reorderBuffer_0_io_loadStoreQueue_2_valid; // @[B4Processor.scala 175:42]
  assign loadStoreQueue_0_io_reorderBuffer_2_bits_destinationTag_threadId = 1'h0; // @[B4Processor.scala 175:42]
  assign loadStoreQueue_0_io_reorderBuffer_2_bits_destinationTag_id =
    reorderBuffer_0_io_loadStoreQueue_2_bits_destinationTag_id; // @[B4Processor.scala 175:42]
  assign loadStoreQueue_0_io_reorderBuffer_3_valid = reorderBuffer_0_io_loadStoreQueue_3_valid; // @[B4Processor.scala 175:42]
  assign loadStoreQueue_0_io_reorderBuffer_3_bits_destinationTag_threadId = 1'h0; // @[B4Processor.scala 175:42]
  assign loadStoreQueue_0_io_reorderBuffer_3_bits_destinationTag_id =
    reorderBuffer_0_io_loadStoreQueue_3_bits_destinationTag_id; // @[B4Processor.scala 175:42]
  assign loadStoreQueue_0_io_memory_ready = dataMemoryBuffer_io_dataIn_0_ready; // @[B4Processor.scala 169:37]
  assign loadStoreQueue_1_clock = clock;
  assign loadStoreQueue_1_reset = reset;
  assign loadStoreQueue_1_io_decoders_0_valid = decoders_1_0_io_loadStoreQueue_valid; // @[B4Processor.scala 149:42]
  assign loadStoreQueue_1_io_decoders_0_bits_accessInfo_accessType =
    decoders_1_0_io_loadStoreQueue_bits_accessInfo_accessType; // @[B4Processor.scala 149:42]
  assign loadStoreQueue_1_io_decoders_0_bits_accessInfo_signed = decoders_1_0_io_loadStoreQueue_bits_accessInfo_signed; // @[B4Processor.scala 149:42]
  assign loadStoreQueue_1_io_decoders_0_bits_accessInfo_accessWidth =
    decoders_1_0_io_loadStoreQueue_bits_accessInfo_accessWidth; // @[B4Processor.scala 149:42]
  assign loadStoreQueue_1_io_decoders_0_bits_addressAndLoadResultTag_threadId =
    decoders_1_0_io_loadStoreQueue_bits_addressAndLoadResultTag_threadId; // @[B4Processor.scala 149:42]
  assign loadStoreQueue_1_io_decoders_0_bits_addressAndLoadResultTag_id =
    decoders_1_0_io_loadStoreQueue_bits_addressAndLoadResultTag_id; // @[B4Processor.scala 149:42]
  assign loadStoreQueue_1_io_decoders_0_bits_address = decoders_1_0_io_loadStoreQueue_bits_address; // @[B4Processor.scala 149:42]
  assign loadStoreQueue_1_io_decoders_0_bits_addressValid = decoders_1_0_io_loadStoreQueue_bits_addressValid; // @[B4Processor.scala 149:42]
  assign loadStoreQueue_1_io_decoders_0_bits_storeDataTag_threadId =
    decoders_1_0_io_loadStoreQueue_bits_storeDataTag_threadId; // @[B4Processor.scala 149:42]
  assign loadStoreQueue_1_io_decoders_0_bits_storeDataTag_id = decoders_1_0_io_loadStoreQueue_bits_storeDataTag_id; // @[B4Processor.scala 149:42]
  assign loadStoreQueue_1_io_decoders_0_bits_storeData = decoders_1_0_io_loadStoreQueue_bits_storeData; // @[B4Processor.scala 149:42]
  assign loadStoreQueue_1_io_decoders_0_bits_storeDataValid = decoders_1_0_io_loadStoreQueue_bits_storeDataValid; // @[B4Processor.scala 149:42]
  assign loadStoreQueue_1_io_outputCollector_outputs_valid = outputCollector_io_outputs_1_outputs_valid; // @[B4Processor.scala 157:44]
  assign loadStoreQueue_1_io_outputCollector_outputs_bits_resultType =
    outputCollector_io_outputs_1_outputs_bits_resultType; // @[B4Processor.scala 157:44]
  assign loadStoreQueue_1_io_outputCollector_outputs_bits_value = outputCollector_io_outputs_1_outputs_bits_value; // @[B4Processor.scala 157:44]
  assign loadStoreQueue_1_io_outputCollector_outputs_bits_tag_threadId =
    outputCollector_io_outputs_1_outputs_bits_tag_threadId; // @[B4Processor.scala 157:44]
  assign loadStoreQueue_1_io_outputCollector_outputs_bits_tag_id = outputCollector_io_outputs_1_outputs_bits_tag_id; // @[B4Processor.scala 157:44]
  assign loadStoreQueue_1_io_reorderBuffer_0_valid = reorderBuffer_1_io_loadStoreQueue_0_valid; // @[B4Processor.scala 175:42]
  assign loadStoreQueue_1_io_reorderBuffer_0_bits_destinationTag_threadId = 1'h1; // @[B4Processor.scala 175:42]
  assign loadStoreQueue_1_io_reorderBuffer_0_bits_destinationTag_id =
    reorderBuffer_1_io_loadStoreQueue_0_bits_destinationTag_id; // @[B4Processor.scala 175:42]
  assign loadStoreQueue_1_io_reorderBuffer_1_valid = reorderBuffer_1_io_loadStoreQueue_1_valid; // @[B4Processor.scala 175:42]
  assign loadStoreQueue_1_io_reorderBuffer_1_bits_destinationTag_threadId = 1'h1; // @[B4Processor.scala 175:42]
  assign loadStoreQueue_1_io_reorderBuffer_1_bits_destinationTag_id =
    reorderBuffer_1_io_loadStoreQueue_1_bits_destinationTag_id; // @[B4Processor.scala 175:42]
  assign loadStoreQueue_1_io_reorderBuffer_2_valid = reorderBuffer_1_io_loadStoreQueue_2_valid; // @[B4Processor.scala 175:42]
  assign loadStoreQueue_1_io_reorderBuffer_2_bits_destinationTag_threadId = 1'h1; // @[B4Processor.scala 175:42]
  assign loadStoreQueue_1_io_reorderBuffer_2_bits_destinationTag_id =
    reorderBuffer_1_io_loadStoreQueue_2_bits_destinationTag_id; // @[B4Processor.scala 175:42]
  assign loadStoreQueue_1_io_reorderBuffer_3_valid = reorderBuffer_1_io_loadStoreQueue_3_valid; // @[B4Processor.scala 175:42]
  assign loadStoreQueue_1_io_reorderBuffer_3_bits_destinationTag_threadId = 1'h1; // @[B4Processor.scala 175:42]
  assign loadStoreQueue_1_io_reorderBuffer_3_bits_destinationTag_id =
    reorderBuffer_1_io_loadStoreQueue_3_bits_destinationTag_id; // @[B4Processor.scala 175:42]
  assign loadStoreQueue_1_io_memory_ready = dataMemoryBuffer_io_dataIn_1_ready; // @[B4Processor.scala 169:37]
  assign dataMemoryBuffer_clock = clock;
  assign dataMemoryBuffer_reset = reset;
  assign dataMemoryBuffer_io_dataIn_0_valid = loadStoreQueue_0_io_memory_valid; // @[B4Processor.scala 169:37]
  assign dataMemoryBuffer_io_dataIn_0_bits_address = loadStoreQueue_0_io_memory_bits_address; // @[B4Processor.scala 169:37]
  assign dataMemoryBuffer_io_dataIn_0_bits_tag_threadId = loadStoreQueue_0_io_memory_bits_tag_threadId; // @[B4Processor.scala 169:37]
  assign dataMemoryBuffer_io_dataIn_0_bits_tag_id = loadStoreQueue_0_io_memory_bits_tag_id; // @[B4Processor.scala 169:37]
  assign dataMemoryBuffer_io_dataIn_0_bits_data = loadStoreQueue_0_io_memory_bits_data; // @[B4Processor.scala 169:37]
  assign dataMemoryBuffer_io_dataIn_0_bits_accessInfo_accessType = loadStoreQueue_0_io_memory_bits_accessInfo_accessType
    ; // @[B4Processor.scala 169:37]
  assign dataMemoryBuffer_io_dataIn_0_bits_accessInfo_signed = loadStoreQueue_0_io_memory_bits_accessInfo_signed; // @[B4Processor.scala 169:37]
  assign dataMemoryBuffer_io_dataIn_0_bits_accessInfo_accessWidth =
    loadStoreQueue_0_io_memory_bits_accessInfo_accessWidth; // @[B4Processor.scala 169:37]
  assign dataMemoryBuffer_io_dataIn_1_valid = loadStoreQueue_1_io_memory_valid; // @[B4Processor.scala 169:37]
  assign dataMemoryBuffer_io_dataIn_1_bits_address = loadStoreQueue_1_io_memory_bits_address; // @[B4Processor.scala 169:37]
  assign dataMemoryBuffer_io_dataIn_1_bits_tag_threadId = loadStoreQueue_1_io_memory_bits_tag_threadId; // @[B4Processor.scala 169:37]
  assign dataMemoryBuffer_io_dataIn_1_bits_tag_id = loadStoreQueue_1_io_memory_bits_tag_id; // @[B4Processor.scala 169:37]
  assign dataMemoryBuffer_io_dataIn_1_bits_data = loadStoreQueue_1_io_memory_bits_data; // @[B4Processor.scala 169:37]
  assign dataMemoryBuffer_io_dataIn_1_bits_accessInfo_accessType = loadStoreQueue_1_io_memory_bits_accessInfo_accessType
    ; // @[B4Processor.scala 169:37]
  assign dataMemoryBuffer_io_dataIn_1_bits_accessInfo_signed = loadStoreQueue_1_io_memory_bits_accessInfo_signed; // @[B4Processor.scala 169:37]
  assign dataMemoryBuffer_io_dataIn_1_bits_accessInfo_accessWidth =
    loadStoreQueue_1_io_memory_bits_accessInfo_accessWidth; // @[B4Processor.scala 169:37]
  assign dataMemoryBuffer_io_dataReadRequest_ready = externalMemoryInterface_io_dataReadRequests_ready; // @[B4Processor.scala 190:47]
  assign dataMemoryBuffer_io_dataWriteRequest_ready = externalMemoryInterface_io_dataWriteRequests_ready; // @[B4Processor.scala 191:48]
  assign outputCollector_clock = clock;
  assign outputCollector_reset = reset;
  assign outputCollector_io_executor_0_valid = executors_0_io_out_valid; // @[B4Processor.scala 89:36]
  assign outputCollector_io_executor_0_bits_resultType = executors_0_io_out_bits_resultType; // @[B4Processor.scala 89:36]
  assign outputCollector_io_executor_0_bits_value = executors_0_io_out_bits_value; // @[B4Processor.scala 89:36]
  assign outputCollector_io_executor_0_bits_tag_threadId = executors_0_io_out_bits_tag_threadId; // @[B4Processor.scala 89:36]
  assign outputCollector_io_executor_0_bits_tag_id = executors_0_io_out_bits_tag_id; // @[B4Processor.scala 89:36]
  assign outputCollector_io_executor_1_valid = executors_1_io_out_valid; // @[B4Processor.scala 89:36]
  assign outputCollector_io_executor_1_bits_resultType = executors_1_io_out_bits_resultType; // @[B4Processor.scala 89:36]
  assign outputCollector_io_executor_1_bits_value = executors_1_io_out_bits_value; // @[B4Processor.scala 89:36]
  assign outputCollector_io_executor_1_bits_tag_threadId = executors_1_io_out_bits_tag_threadId; // @[B4Processor.scala 89:36]
  assign outputCollector_io_executor_1_bits_tag_id = executors_1_io_out_bits_tag_id; // @[B4Processor.scala 89:36]
  assign outputCollector_io_dataMemory_valid = externalMemoryInterface_io_dataReadOut_valid; // @[B4Processor.scala 68:33]
  assign outputCollector_io_dataMemory_bits_value = externalMemoryInterface_io_dataReadOut_bits_value; // @[B4Processor.scala 68:33]
  assign outputCollector_io_dataMemory_bits_isError = externalMemoryInterface_io_dataReadOut_bits_isError; // @[B4Processor.scala 68:33]
  assign outputCollector_io_dataMemory_bits_tag_threadId = externalMemoryInterface_io_dataReadOut_bits_tag_threadId; // @[B4Processor.scala 68:33]
  assign outputCollector_io_dataMemory_bits_tag_id = externalMemoryInterface_io_dataReadOut_bits_tag_id; // @[B4Processor.scala 68:33]
  assign outputCollector_io_csr_0_valid = csr_0_io_CSROutput_valid; // @[B4Processor.scala 108:27]
  assign outputCollector_io_csr_0_bits_value = csr_0_io_CSROutput_bits_value; // @[B4Processor.scala 108:27]
  assign outputCollector_io_csr_0_bits_isError = csr_0_io_CSROutput_bits_isError; // @[B4Processor.scala 108:27]
  assign outputCollector_io_csr_0_bits_tag_threadId = csr_0_io_CSROutput_bits_tag_threadId; // @[B4Processor.scala 108:27]
  assign outputCollector_io_csr_0_bits_tag_id = csr_0_io_CSROutput_bits_tag_id; // @[B4Processor.scala 108:27]
  assign outputCollector_io_csr_1_valid = csr_1_io_CSROutput_valid; // @[B4Processor.scala 108:27]
  assign outputCollector_io_csr_1_bits_value = csr_1_io_CSROutput_bits_value; // @[B4Processor.scala 108:27]
  assign outputCollector_io_csr_1_bits_isError = csr_1_io_CSROutput_bits_isError; // @[B4Processor.scala 108:27]
  assign outputCollector_io_csr_1_bits_tag_threadId = csr_1_io_CSROutput_bits_tag_threadId; // @[B4Processor.scala 108:27]
  assign outputCollector_io_csr_1_bits_tag_id = csr_1_io_CSROutput_bits_tag_id; // @[B4Processor.scala 108:27]
  assign outputCollector_io_isError_0 = reorderBuffer_0_io_isError; // @[B4Processor.scala 119:37]
  assign outputCollector_io_isError_1 = reorderBuffer_1_io_isError; // @[B4Processor.scala 119:37]
  assign branchAddressCollector_clock = clock;
  assign branchAddressCollector_reset = reset;
  assign branchAddressCollector_io_executor_0_valid = executors_0_io_fetch_valid; // @[B4Processor.scala 92:43]
  assign branchAddressCollector_io_executor_0_bits_threadId = executors_0_io_fetch_bits_threadId; // @[B4Processor.scala 92:43]
  assign branchAddressCollector_io_executor_0_bits_programCounterOffset = executors_0_io_fetch_bits_programCounterOffset
    ; // @[B4Processor.scala 92:43]
  assign branchAddressCollector_io_executor_1_valid = executors_1_io_fetch_valid; // @[B4Processor.scala 92:43]
  assign branchAddressCollector_io_executor_1_bits_threadId = executors_1_io_fetch_bits_threadId; // @[B4Processor.scala 92:43]
  assign branchAddressCollector_io_executor_1_bits_programCounterOffset = executors_1_io_fetch_bits_programCounterOffset
    ; // @[B4Processor.scala 92:43]
  assign branchAddressCollector_io_isError_0 = reorderBuffer_0_io_isError; // @[B4Processor.scala 120:44]
  assign branchAddressCollector_io_isError_1 = reorderBuffer_1_io_isError; // @[B4Processor.scala 120:44]
  assign uncompresser_0_0_io_fetch_valid = fetchBuffer_0_io_output_0_valid; // @[B4Processor.scala 127:37]
  assign uncompresser_0_0_io_fetch_bits_instruction = fetchBuffer_0_io_output_0_bits_instruction; // @[B4Processor.scala 127:37]
  assign uncompresser_0_0_io_fetch_bits_programCounter = fetchBuffer_0_io_output_0_bits_programCounter; // @[B4Processor.scala 127:37]
  assign uncompresser_0_0_io_decoder_ready = decoders_0_0_io_instructionFetch_ready; // @[B4Processor.scala 130:44]
  assign uncompresser_1_0_io_fetch_valid = fetchBuffer_1_io_output_0_valid; // @[B4Processor.scala 127:37]
  assign uncompresser_1_0_io_fetch_bits_instruction = fetchBuffer_1_io_output_0_bits_instruction; // @[B4Processor.scala 127:37]
  assign uncompresser_1_0_io_fetch_bits_programCounter = fetchBuffer_1_io_output_0_bits_programCounter; // @[B4Processor.scala 127:37]
  assign uncompresser_1_0_io_decoder_ready = decoders_1_0_io_instructionFetch_ready; // @[B4Processor.scala 130:44]
  assign decoders_0_0_io_instructionFetch_valid = uncompresser_0_0_io_decoder_valid; // @[B4Processor.scala 130:44]
  assign decoders_0_0_io_instructionFetch_bits_instruction = uncompresser_0_0_io_decoder_bits_instruction; // @[B4Processor.scala 130:44]
  assign decoders_0_0_io_instructionFetch_bits_programCounter = uncompresser_0_0_io_decoder_bits_programCounter; // @[B4Processor.scala 130:44]
  assign decoders_0_0_io_instructionFetch_bits_wasCompressed = uncompresser_0_0_io_decoder_bits_wasCompressed; // @[B4Processor.scala 130:44]
  assign decoders_0_0_io_reorderBuffer_source1_matchingTag_valid =
    reorderBuffer_0_io_decoders_0_source1_matchingTag_valid; // @[B4Processor.scala 133:41]
  assign decoders_0_0_io_reorderBuffer_source1_matchingTag_bits_id =
    reorderBuffer_0_io_decoders_0_source1_matchingTag_bits_id; // @[B4Processor.scala 133:41]
  assign decoders_0_0_io_reorderBuffer_source1_value_valid = reorderBuffer_0_io_decoders_0_source1_value_valid; // @[B4Processor.scala 133:41]
  assign decoders_0_0_io_reorderBuffer_source1_value_bits = reorderBuffer_0_io_decoders_0_source1_value_bits; // @[B4Processor.scala 133:41]
  assign decoders_0_0_io_reorderBuffer_source2_matchingTag_valid =
    reorderBuffer_0_io_decoders_0_source2_matchingTag_valid; // @[B4Processor.scala 133:41]
  assign decoders_0_0_io_reorderBuffer_source2_matchingTag_bits_id =
    reorderBuffer_0_io_decoders_0_source2_matchingTag_bits_id; // @[B4Processor.scala 133:41]
  assign decoders_0_0_io_reorderBuffer_source2_value_valid = reorderBuffer_0_io_decoders_0_source2_value_valid; // @[B4Processor.scala 133:41]
  assign decoders_0_0_io_reorderBuffer_source2_value_bits = reorderBuffer_0_io_decoders_0_source2_value_bits; // @[B4Processor.scala 133:41]
  assign decoders_0_0_io_reorderBuffer_destination_destinationTag_id =
    reorderBuffer_0_io_decoders_0_destination_destinationTag_id; // @[B4Processor.scala 133:41]
  assign decoders_0_0_io_reorderBuffer_ready = reorderBuffer_0_io_decoders_0_ready; // @[B4Processor.scala 133:41]
  assign decoders_0_0_io_outputCollector_outputs_valid = outputCollector_io_outputs_0_outputs_valid; // @[B4Processor.scala 146:43]
  assign decoders_0_0_io_outputCollector_outputs_bits_resultType = outputCollector_io_outputs_0_outputs_bits_resultType; // @[B4Processor.scala 146:43]
  assign decoders_0_0_io_outputCollector_outputs_bits_value = outputCollector_io_outputs_0_outputs_bits_value; // @[B4Processor.scala 146:43]
  assign decoders_0_0_io_outputCollector_outputs_bits_tag_threadId =
    outputCollector_io_outputs_0_outputs_bits_tag_threadId; // @[B4Processor.scala 146:43]
  assign decoders_0_0_io_outputCollector_outputs_bits_tag_id = outputCollector_io_outputs_0_outputs_bits_tag_id; // @[B4Processor.scala 146:43]
  assign decoders_0_0_io_registerFile_value1 = registerFile_0_io_decoders_0_value1; // @[B4Processor.scala 140:40]
  assign decoders_0_0_io_registerFile_value2 = registerFile_0_io_decoders_0_value2; // @[B4Processor.scala 140:40]
  assign decoders_0_0_io_reservationStation_ready = reservationStation_io_decoder_0_ready; // @[B4Processor.scala 136:46]
  assign decoders_0_0_io_loadStoreQueue_ready = loadStoreQueue_0_io_decoders_0_ready; // @[B4Processor.scala 149:42]
  assign decoders_0_0_io_csr_ready = csrReservationStation_0_io_decoderInput_0_ready; // @[B4Processor.scala 125:31]
  assign decoders_1_0_io_instructionFetch_valid = uncompresser_1_0_io_decoder_valid; // @[B4Processor.scala 130:44]
  assign decoders_1_0_io_instructionFetch_bits_instruction = uncompresser_1_0_io_decoder_bits_instruction; // @[B4Processor.scala 130:44]
  assign decoders_1_0_io_instructionFetch_bits_programCounter = uncompresser_1_0_io_decoder_bits_programCounter; // @[B4Processor.scala 130:44]
  assign decoders_1_0_io_instructionFetch_bits_wasCompressed = uncompresser_1_0_io_decoder_bits_wasCompressed; // @[B4Processor.scala 130:44]
  assign decoders_1_0_io_reorderBuffer_source1_matchingTag_valid =
    reorderBuffer_1_io_decoders_0_source1_matchingTag_valid; // @[B4Processor.scala 133:41]
  assign decoders_1_0_io_reorderBuffer_source1_matchingTag_bits_id =
    reorderBuffer_1_io_decoders_0_source1_matchingTag_bits_id; // @[B4Processor.scala 133:41]
  assign decoders_1_0_io_reorderBuffer_source1_value_valid = reorderBuffer_1_io_decoders_0_source1_value_valid; // @[B4Processor.scala 133:41]
  assign decoders_1_0_io_reorderBuffer_source1_value_bits = reorderBuffer_1_io_decoders_0_source1_value_bits; // @[B4Processor.scala 133:41]
  assign decoders_1_0_io_reorderBuffer_source2_matchingTag_valid =
    reorderBuffer_1_io_decoders_0_source2_matchingTag_valid; // @[B4Processor.scala 133:41]
  assign decoders_1_0_io_reorderBuffer_source2_matchingTag_bits_id =
    reorderBuffer_1_io_decoders_0_source2_matchingTag_bits_id; // @[B4Processor.scala 133:41]
  assign decoders_1_0_io_reorderBuffer_source2_value_valid = reorderBuffer_1_io_decoders_0_source2_value_valid; // @[B4Processor.scala 133:41]
  assign decoders_1_0_io_reorderBuffer_source2_value_bits = reorderBuffer_1_io_decoders_0_source2_value_bits; // @[B4Processor.scala 133:41]
  assign decoders_1_0_io_reorderBuffer_destination_destinationTag_id =
    reorderBuffer_1_io_decoders_0_destination_destinationTag_id; // @[B4Processor.scala 133:41]
  assign decoders_1_0_io_reorderBuffer_ready = reorderBuffer_1_io_decoders_0_ready; // @[B4Processor.scala 133:41]
  assign decoders_1_0_io_outputCollector_outputs_valid = outputCollector_io_outputs_1_outputs_valid; // @[B4Processor.scala 146:43]
  assign decoders_1_0_io_outputCollector_outputs_bits_resultType = outputCollector_io_outputs_1_outputs_bits_resultType; // @[B4Processor.scala 146:43]
  assign decoders_1_0_io_outputCollector_outputs_bits_value = outputCollector_io_outputs_1_outputs_bits_value; // @[B4Processor.scala 146:43]
  assign decoders_1_0_io_outputCollector_outputs_bits_tag_threadId =
    outputCollector_io_outputs_1_outputs_bits_tag_threadId; // @[B4Processor.scala 146:43]
  assign decoders_1_0_io_outputCollector_outputs_bits_tag_id = outputCollector_io_outputs_1_outputs_bits_tag_id; // @[B4Processor.scala 146:43]
  assign decoders_1_0_io_registerFile_value1 = registerFile_1_io_decoders_0_value1; // @[B4Processor.scala 140:40]
  assign decoders_1_0_io_registerFile_value2 = registerFile_1_io_decoders_0_value2; // @[B4Processor.scala 140:40]
  assign decoders_1_0_io_reservationStation_ready = reservationStation_io_decoder_1_ready; // @[B4Processor.scala 136:46]
  assign decoders_1_0_io_loadStoreQueue_ready = loadStoreQueue_1_io_decoders_0_ready; // @[B4Processor.scala 149:42]
  assign decoders_1_0_io_csr_ready = csrReservationStation_1_io_decoderInput_0_ready; // @[B4Processor.scala 125:31]
  assign reservationStation_clock = clock;
  assign reservationStation_reset = reset;
  assign reservationStation_io_collectedOutput_0_outputs_valid = outputCollector_io_outputs_0_outputs_valid; // @[B4Processor.scala 96:41]
  assign reservationStation_io_collectedOutput_0_outputs_bits_resultType =
    outputCollector_io_outputs_0_outputs_bits_resultType; // @[B4Processor.scala 96:41]
  assign reservationStation_io_collectedOutput_0_outputs_bits_value = outputCollector_io_outputs_0_outputs_bits_value; // @[B4Processor.scala 96:41]
  assign reservationStation_io_collectedOutput_0_outputs_bits_tag_threadId =
    outputCollector_io_outputs_0_outputs_bits_tag_threadId; // @[B4Processor.scala 96:41]
  assign reservationStation_io_collectedOutput_0_outputs_bits_tag_id = outputCollector_io_outputs_0_outputs_bits_tag_id; // @[B4Processor.scala 96:41]
  assign reservationStation_io_collectedOutput_1_outputs_valid = outputCollector_io_outputs_1_outputs_valid; // @[B4Processor.scala 96:41]
  assign reservationStation_io_collectedOutput_1_outputs_bits_resultType =
    outputCollector_io_outputs_1_outputs_bits_resultType; // @[B4Processor.scala 96:41]
  assign reservationStation_io_collectedOutput_1_outputs_bits_value = outputCollector_io_outputs_1_outputs_bits_value; // @[B4Processor.scala 96:41]
  assign reservationStation_io_collectedOutput_1_outputs_bits_tag_threadId =
    outputCollector_io_outputs_1_outputs_bits_tag_threadId; // @[B4Processor.scala 96:41]
  assign reservationStation_io_collectedOutput_1_outputs_bits_tag_id = outputCollector_io_outputs_1_outputs_bits_tag_id; // @[B4Processor.scala 96:41]
  assign reservationStation_io_executor_0_ready = executors_0_io_reservationStation_ready; // @[B4Processor.scala 86:39]
  assign reservationStation_io_executor_1_ready = executors_1_io_reservationStation_ready; // @[B4Processor.scala 86:39]
  assign reservationStation_io_decoder_0_entry_opcode = decoders_0_0_io_reservationStation_entry_opcode; // @[B4Processor.scala 136:46]
  assign reservationStation_io_decoder_0_entry_function3 = decoders_0_0_io_reservationStation_entry_function3; // @[B4Processor.scala 136:46]
  assign reservationStation_io_decoder_0_entry_immediateOrFunction7 =
    decoders_0_0_io_reservationStation_entry_immediateOrFunction7; // @[B4Processor.scala 136:46]
  assign reservationStation_io_decoder_0_entry_sourceTag1_threadId =
    decoders_0_0_io_reservationStation_entry_sourceTag1_threadId; // @[B4Processor.scala 136:46]
  assign reservationStation_io_decoder_0_entry_sourceTag1_id = decoders_0_0_io_reservationStation_entry_sourceTag1_id; // @[B4Processor.scala 136:46]
  assign reservationStation_io_decoder_0_entry_ready1 = decoders_0_0_io_reservationStation_entry_ready1; // @[B4Processor.scala 136:46]
  assign reservationStation_io_decoder_0_entry_value1 = decoders_0_0_io_reservationStation_entry_value1; // @[B4Processor.scala 136:46]
  assign reservationStation_io_decoder_0_entry_sourceTag2_threadId =
    decoders_0_0_io_reservationStation_entry_sourceTag2_threadId; // @[B4Processor.scala 136:46]
  assign reservationStation_io_decoder_0_entry_sourceTag2_id = decoders_0_0_io_reservationStation_entry_sourceTag2_id; // @[B4Processor.scala 136:46]
  assign reservationStation_io_decoder_0_entry_ready2 = decoders_0_0_io_reservationStation_entry_ready2; // @[B4Processor.scala 136:46]
  assign reservationStation_io_decoder_0_entry_value2 = decoders_0_0_io_reservationStation_entry_value2; // @[B4Processor.scala 136:46]
  assign reservationStation_io_decoder_0_entry_destinationTag_id =
    decoders_0_0_io_reservationStation_entry_destinationTag_id; // @[B4Processor.scala 136:46]
  assign reservationStation_io_decoder_0_entry_wasCompressed = decoders_0_0_io_reservationStation_entry_wasCompressed; // @[B4Processor.scala 136:46]
  assign reservationStation_io_decoder_0_entry_valid = decoders_0_0_io_reservationStation_entry_valid; // @[B4Processor.scala 136:46]
  assign reservationStation_io_decoder_1_entry_opcode = decoders_1_0_io_reservationStation_entry_opcode; // @[B4Processor.scala 136:46]
  assign reservationStation_io_decoder_1_entry_function3 = decoders_1_0_io_reservationStation_entry_function3; // @[B4Processor.scala 136:46]
  assign reservationStation_io_decoder_1_entry_immediateOrFunction7 =
    decoders_1_0_io_reservationStation_entry_immediateOrFunction7; // @[B4Processor.scala 136:46]
  assign reservationStation_io_decoder_1_entry_sourceTag1_threadId =
    decoders_1_0_io_reservationStation_entry_sourceTag1_threadId; // @[B4Processor.scala 136:46]
  assign reservationStation_io_decoder_1_entry_sourceTag1_id = decoders_1_0_io_reservationStation_entry_sourceTag1_id; // @[B4Processor.scala 136:46]
  assign reservationStation_io_decoder_1_entry_ready1 = decoders_1_0_io_reservationStation_entry_ready1; // @[B4Processor.scala 136:46]
  assign reservationStation_io_decoder_1_entry_value1 = decoders_1_0_io_reservationStation_entry_value1; // @[B4Processor.scala 136:46]
  assign reservationStation_io_decoder_1_entry_sourceTag2_threadId =
    decoders_1_0_io_reservationStation_entry_sourceTag2_threadId; // @[B4Processor.scala 136:46]
  assign reservationStation_io_decoder_1_entry_sourceTag2_id = decoders_1_0_io_reservationStation_entry_sourceTag2_id; // @[B4Processor.scala 136:46]
  assign reservationStation_io_decoder_1_entry_ready2 = decoders_1_0_io_reservationStation_entry_ready2; // @[B4Processor.scala 136:46]
  assign reservationStation_io_decoder_1_entry_value2 = decoders_1_0_io_reservationStation_entry_value2; // @[B4Processor.scala 136:46]
  assign reservationStation_io_decoder_1_entry_destinationTag_id =
    decoders_1_0_io_reservationStation_entry_destinationTag_id; // @[B4Processor.scala 136:46]
  assign reservationStation_io_decoder_1_entry_wasCompressed = decoders_1_0_io_reservationStation_entry_wasCompressed; // @[B4Processor.scala 136:46]
  assign reservationStation_io_decoder_1_entry_valid = decoders_1_0_io_reservationStation_entry_valid; // @[B4Processor.scala 136:46]
  assign executors_0_io_reservationStation_valid = reservationStation_io_executor_0_valid; // @[B4Processor.scala 86:39]
  assign executors_0_io_reservationStation_bits_destinationTag_threadId =
    reservationStation_io_executor_0_bits_destinationTag_threadId; // @[B4Processor.scala 86:39]
  assign executors_0_io_reservationStation_bits_destinationTag_id =
    reservationStation_io_executor_0_bits_destinationTag_id; // @[B4Processor.scala 86:39]
  assign executors_0_io_reservationStation_bits_value1 = reservationStation_io_executor_0_bits_value1; // @[B4Processor.scala 86:39]
  assign executors_0_io_reservationStation_bits_value2 = reservationStation_io_executor_0_bits_value2; // @[B4Processor.scala 86:39]
  assign executors_0_io_reservationStation_bits_function3 = reservationStation_io_executor_0_bits_function3; // @[B4Processor.scala 86:39]
  assign executors_0_io_reservationStation_bits_immediateOrFunction7 =
    reservationStation_io_executor_0_bits_immediateOrFunction7; // @[B4Processor.scala 86:39]
  assign executors_0_io_reservationStation_bits_opcode = reservationStation_io_executor_0_bits_opcode; // @[B4Processor.scala 86:39]
  assign executors_0_io_reservationStation_bits_wasCompressed = reservationStation_io_executor_0_bits_wasCompressed; // @[B4Processor.scala 86:39]
  assign executors_0_io_out_ready = outputCollector_io_executor_0_ready; // @[B4Processor.scala 89:36]
  assign executors_0_io_fetch_ready = branchAddressCollector_io_executor_0_ready; // @[B4Processor.scala 92:43]
  assign executors_1_io_reservationStation_valid = reservationStation_io_executor_1_valid; // @[B4Processor.scala 86:39]
  assign executors_1_io_reservationStation_bits_destinationTag_threadId =
    reservationStation_io_executor_1_bits_destinationTag_threadId; // @[B4Processor.scala 86:39]
  assign executors_1_io_reservationStation_bits_destinationTag_id =
    reservationStation_io_executor_1_bits_destinationTag_id; // @[B4Processor.scala 86:39]
  assign executors_1_io_reservationStation_bits_value1 = reservationStation_io_executor_1_bits_value1; // @[B4Processor.scala 86:39]
  assign executors_1_io_reservationStation_bits_value2 = reservationStation_io_executor_1_bits_value2; // @[B4Processor.scala 86:39]
  assign executors_1_io_reservationStation_bits_function3 = reservationStation_io_executor_1_bits_function3; // @[B4Processor.scala 86:39]
  assign executors_1_io_reservationStation_bits_immediateOrFunction7 =
    reservationStation_io_executor_1_bits_immediateOrFunction7; // @[B4Processor.scala 86:39]
  assign executors_1_io_reservationStation_bits_opcode = reservationStation_io_executor_1_bits_opcode; // @[B4Processor.scala 86:39]
  assign executors_1_io_reservationStation_bits_wasCompressed = reservationStation_io_executor_1_bits_wasCompressed; // @[B4Processor.scala 86:39]
  assign executors_1_io_out_ready = outputCollector_io_executor_1_ready; // @[B4Processor.scala 89:36]
  assign executors_1_io_fetch_ready = branchAddressCollector_io_executor_1_ready; // @[B4Processor.scala 92:43]
  assign externalMemoryInterface_clock = clock;
  assign externalMemoryInterface_reset = reset;
  assign externalMemoryInterface_io_dataWriteRequests_valid = dataMemoryBuffer_io_dataWriteRequest_valid; // @[B4Processor.scala 191:48]
  assign externalMemoryInterface_io_dataWriteRequests_bits_address = dataMemoryBuffer_io_dataWriteRequest_bits_address; // @[B4Processor.scala 191:48]
  assign externalMemoryInterface_io_dataWriteRequests_bits_data = dataMemoryBuffer_io_dataWriteRequest_bits_data; // @[B4Processor.scala 191:48]
  assign externalMemoryInterface_io_dataWriteRequests_bits_mask = dataMemoryBuffer_io_dataWriteRequest_bits_mask; // @[B4Processor.scala 191:48]
  assign externalMemoryInterface_io_dataReadRequests_valid = dataMemoryBuffer_io_dataReadRequest_valid; // @[B4Processor.scala 190:47]
  assign externalMemoryInterface_io_dataReadRequests_bits_address = dataMemoryBuffer_io_dataReadRequest_bits_address; // @[B4Processor.scala 190:47]
  assign externalMemoryInterface_io_dataReadRequests_bits_size = dataMemoryBuffer_io_dataReadRequest_bits_size; // @[B4Processor.scala 190:47]
  assign externalMemoryInterface_io_dataReadRequests_bits_signed = dataMemoryBuffer_io_dataReadRequest_bits_signed; // @[B4Processor.scala 190:47]
  assign externalMemoryInterface_io_dataReadRequests_bits_outputTag_threadId =
    dataMemoryBuffer_io_dataReadRequest_bits_outputTag_threadId; // @[B4Processor.scala 190:47]
  assign externalMemoryInterface_io_dataReadRequests_bits_outputTag_id =
    dataMemoryBuffer_io_dataReadRequest_bits_outputTag_id; // @[B4Processor.scala 190:47]
  assign externalMemoryInterface_io_instructionFetchRequest_0_valid = instructionCache_0_io_memory_request_valid; // @[B4Processor.scala 178:61]
  assign externalMemoryInterface_io_instructionFetchRequest_0_bits_address =
    instructionCache_0_io_memory_request_bits_address; // @[B4Processor.scala 178:61]
  assign externalMemoryInterface_io_instructionFetchRequest_1_valid = instructionCache_1_io_memory_request_valid; // @[B4Processor.scala 178:61]
  assign externalMemoryInterface_io_instructionFetchRequest_1_bits_address =
    instructionCache_1_io_memory_request_bits_address; // @[B4Processor.scala 178:61]
  assign externalMemoryInterface_io_dataReadOut_ready = outputCollector_io_dataMemory_ready; // @[B4Processor.scala 68:33]
  assign externalMemoryInterface_io_coordinator_writeAddress_ready = axi_writeAddress_ready; // @[B4Processor.scala 65:7]
  assign externalMemoryInterface_io_coordinator_write_ready = axi_write_ready; // @[B4Processor.scala 65:7]
  assign externalMemoryInterface_io_coordinator_writeResponse_valid = axi_writeResponse_valid; // @[B4Processor.scala 65:7]
  assign externalMemoryInterface_io_coordinator_readAddress_ready = axi_readAddress_ready; // @[B4Processor.scala 65:7]
  assign externalMemoryInterface_io_coordinator_read_valid = axi_read_valid; // @[B4Processor.scala 65:7]
  assign externalMemoryInterface_io_coordinator_read_bits_DATA = axi_read_bits_DATA; // @[B4Processor.scala 65:7]
  assign externalMemoryInterface_io_coordinator_read_bits_RESP = axi_read_bits_RESP; // @[B4Processor.scala 65:7]
  assign csrReservationStation_0_clock = clock;
  assign csrReservationStation_0_reset = reset;
  assign csrReservationStation_0_io_decoderInput_0_valid = decoders_0_0_io_csr_valid; // @[B4Processor.scala 125:31]
  assign csrReservationStation_0_io_decoderInput_0_bits_sourceTag_threadId = decoders_0_0_io_csr_bits_sourceTag_threadId
    ; // @[B4Processor.scala 125:31]
  assign csrReservationStation_0_io_decoderInput_0_bits_sourceTag_id = decoders_0_0_io_csr_bits_sourceTag_id; // @[B4Processor.scala 125:31]
  assign csrReservationStation_0_io_decoderInput_0_bits_destinationTag_threadId = 1'h0; // @[B4Processor.scala 125:31]
  assign csrReservationStation_0_io_decoderInput_0_bits_destinationTag_id = decoders_0_0_io_csr_bits_destinationTag_id; // @[B4Processor.scala 125:31]
  assign csrReservationStation_0_io_decoderInput_0_bits_value = decoders_0_0_io_csr_bits_value; // @[B4Processor.scala 125:31]
  assign csrReservationStation_0_io_decoderInput_0_bits_ready = decoders_0_0_io_csr_bits_ready; // @[B4Processor.scala 125:31]
  assign csrReservationStation_0_io_decoderInput_0_bits_address = decoders_0_0_io_csr_bits_address; // @[B4Processor.scala 125:31]
  assign csrReservationStation_0_io_decoderInput_0_bits_csrAccessType = decoders_0_0_io_csr_bits_csrAccessType; // @[B4Processor.scala 125:31]
  assign csrReservationStation_0_io_toCSR_ready = csr_0_io_decoderInput_ready; // @[B4Processor.scala 106:41]
  assign csrReservationStation_0_io_output_outputs_valid = outputCollector_io_outputs_0_outputs_valid; // @[B4Processor.scala 110:42]
  assign csrReservationStation_0_io_output_outputs_bits_value = outputCollector_io_outputs_0_outputs_bits_value; // @[B4Processor.scala 110:42]
  assign csrReservationStation_0_io_output_outputs_bits_tag_threadId =
    outputCollector_io_outputs_0_outputs_bits_tag_threadId; // @[B4Processor.scala 110:42]
  assign csrReservationStation_0_io_output_outputs_bits_tag_id = outputCollector_io_outputs_0_outputs_bits_tag_id; // @[B4Processor.scala 110:42]
  assign csrReservationStation_1_clock = clock;
  assign csrReservationStation_1_reset = reset;
  assign csrReservationStation_1_io_decoderInput_0_valid = decoders_1_0_io_csr_valid; // @[B4Processor.scala 125:31]
  assign csrReservationStation_1_io_decoderInput_0_bits_sourceTag_threadId = decoders_1_0_io_csr_bits_sourceTag_threadId
    ; // @[B4Processor.scala 125:31]
  assign csrReservationStation_1_io_decoderInput_0_bits_sourceTag_id = decoders_1_0_io_csr_bits_sourceTag_id; // @[B4Processor.scala 125:31]
  assign csrReservationStation_1_io_decoderInput_0_bits_destinationTag_threadId = 1'h1; // @[B4Processor.scala 125:31]
  assign csrReservationStation_1_io_decoderInput_0_bits_destinationTag_id = decoders_1_0_io_csr_bits_destinationTag_id; // @[B4Processor.scala 125:31]
  assign csrReservationStation_1_io_decoderInput_0_bits_value = decoders_1_0_io_csr_bits_value; // @[B4Processor.scala 125:31]
  assign csrReservationStation_1_io_decoderInput_0_bits_ready = decoders_1_0_io_csr_bits_ready; // @[B4Processor.scala 125:31]
  assign csrReservationStation_1_io_decoderInput_0_bits_address = decoders_1_0_io_csr_bits_address; // @[B4Processor.scala 125:31]
  assign csrReservationStation_1_io_decoderInput_0_bits_csrAccessType = decoders_1_0_io_csr_bits_csrAccessType; // @[B4Processor.scala 125:31]
  assign csrReservationStation_1_io_toCSR_ready = csr_1_io_decoderInput_ready; // @[B4Processor.scala 106:41]
  assign csrReservationStation_1_io_output_outputs_valid = outputCollector_io_outputs_1_outputs_valid; // @[B4Processor.scala 110:42]
  assign csrReservationStation_1_io_output_outputs_bits_value = outputCollector_io_outputs_1_outputs_bits_value; // @[B4Processor.scala 110:42]
  assign csrReservationStation_1_io_output_outputs_bits_tag_threadId =
    outputCollector_io_outputs_1_outputs_bits_tag_threadId; // @[B4Processor.scala 110:42]
  assign csrReservationStation_1_io_output_outputs_bits_tag_id = outputCollector_io_outputs_1_outputs_bits_tag_id; // @[B4Processor.scala 110:42]
  assign csr_0_clock = clock;
  assign csr_0_reset = reset;
  assign csr_0_io_decoderInput_valid = csrReservationStation_0_io_toCSR_valid; // @[B4Processor.scala 106:41]
  assign csr_0_io_decoderInput_bits_address = csrReservationStation_0_io_toCSR_bits_address; // @[B4Processor.scala 106:41]
  assign csr_0_io_decoderInput_bits_value = csrReservationStation_0_io_toCSR_bits_value; // @[B4Processor.scala 106:41]
  assign csr_0_io_decoderInput_bits_destinationTag_threadId =
    csrReservationStation_0_io_toCSR_bits_destinationTag_threadId; // @[B4Processor.scala 106:41]
  assign csr_0_io_decoderInput_bits_destinationTag_id = csrReservationStation_0_io_toCSR_bits_destinationTag_id; // @[B4Processor.scala 106:41]
  assign csr_0_io_decoderInput_bits_csrAccessType = csrReservationStation_0_io_toCSR_bits_csrAccessType; // @[B4Processor.scala 106:41]
  assign csr_0_io_CSROutput_ready = outputCollector_io_csr_0_ready; // @[B4Processor.scala 108:27]
  assign csr_0_io_reorderBuffer_retireCount = reorderBuffer_0_io_csr_retireCount; // @[B4Processor.scala 112:31]
  assign csr_1_clock = clock;
  assign csr_1_reset = reset;
  assign csr_1_io_decoderInput_valid = csrReservationStation_1_io_toCSR_valid; // @[B4Processor.scala 106:41]
  assign csr_1_io_decoderInput_bits_address = csrReservationStation_1_io_toCSR_bits_address; // @[B4Processor.scala 106:41]
  assign csr_1_io_decoderInput_bits_value = csrReservationStation_1_io_toCSR_bits_value; // @[B4Processor.scala 106:41]
  assign csr_1_io_decoderInput_bits_destinationTag_threadId =
    csrReservationStation_1_io_toCSR_bits_destinationTag_threadId; // @[B4Processor.scala 106:41]
  assign csr_1_io_decoderInput_bits_destinationTag_id = csrReservationStation_1_io_toCSR_bits_destinationTag_id; // @[B4Processor.scala 106:41]
  assign csr_1_io_decoderInput_bits_csrAccessType = csrReservationStation_1_io_toCSR_bits_csrAccessType; // @[B4Processor.scala 106:41]
  assign csr_1_io_CSROutput_ready = outputCollector_io_csr_1_ready; // @[B4Processor.scala 108:27]
  assign csr_1_io_reorderBuffer_retireCount = reorderBuffer_1_io_csr_retireCount; // @[B4Processor.scala 112:31]
endmodule
